// Generated using mul32_gen.swift

`timescale 1ns/1ns

module ArrayMultiplier(A, B, Z);

input [31: 0] A, B;
output [63: 0] Z;

wire [31:0] sum0;
wire [31:0] sum1;
wire [31:0] sum2;
wire [31:0] sum3;
wire [31:0] sum4;
wire [31:0] sum5;
wire [31:0] sum6;
wire [31:0] sum7;
wire [31:0] sum8;
wire [31:0] sum9;
wire [31:0] sum10;
wire [31:0] sum11;
wire [31:0] sum12;
wire [31:0] sum13;
wire [31:0] sum14;
wire [31:0] sum15;
wire [31:0] sum16;
wire [31:0] sum17;
wire [31:0] sum18;
wire [31:0] sum19;
wire [31:0] sum20;
wire [31:0] sum21;
wire [31:0] sum22;
wire [31:0] sum23;
wire [31:0] sum24;
wire [31:0] sum25;
wire [31:0] sum26;
wire [31:0] sum27;
wire [31:0] sum28;
wire [31:0] sum29;
wire [31:0] sum30;
wire [31:0] sum31;
assign sum0 = A & {32{B[0]}};

wire [31:0] carry0;
wire [31:0] carry1;
wire [31:0] carry2;
wire [31:0] carry3;
wire [31:0] carry4;
wire [31:0] carry5;
wire [31:0] carry6;
wire [31:0] carry7;
wire [31:0] carry8;
wire [31:0] carry9;
wire [31:0] carry10;
wire [31:0] carry11;
wire [31:0] carry12;
wire [31:0] carry13;
wire [31:0] carry14;
wire [31:0] carry15;
wire [31:0] carry16;
wire [31:0] carry17;
wire [31:0] carry18;
wire [31:0] carry19;
wire [31:0] carry20;
wire [31:0] carry21;
wire [31:0] carry22;
wire [31:0] carry23;
wire [31:0] carry24;
wire [31:0] carry25;
wire [31:0] carry26;
wire [31:0] carry27;
wire [31:0] carry28;
wire [31:0] carry29;
wire [31:0] carry30;
wire [31:0] carry31;
assign carry0 = 32'b0;

FA fa1_0(.a(sum0[1]), .b(A[0] & B[1]), .ci(1'b0), .s(Z[1]), .co(carry1[0]));
FA fa1_1(.a(sum0[2]), .b(A[1] & B[1]), .ci(carry1[0]), .s(sum1[1]), .co(carry1[1]));
FA fa1_2(.a(sum0[3]), .b(A[2] & B[1]), .ci(carry1[1]), .s(sum1[2]), .co(carry1[2]));
FA fa1_3(.a(sum0[4]), .b(A[3] & B[1]), .ci(carry1[2]), .s(sum1[3]), .co(carry1[3]));
FA fa1_4(.a(sum0[5]), .b(A[4] & B[1]), .ci(carry1[3]), .s(sum1[4]), .co(carry1[4]));
FA fa1_5(.a(sum0[6]), .b(A[5] & B[1]), .ci(carry1[4]), .s(sum1[5]), .co(carry1[5]));
FA fa1_6(.a(sum0[7]), .b(A[6] & B[1]), .ci(carry1[5]), .s(sum1[6]), .co(carry1[6]));
FA fa1_7(.a(sum0[8]), .b(A[7] & B[1]), .ci(carry1[6]), .s(sum1[7]), .co(carry1[7]));
FA fa1_8(.a(sum0[9]), .b(A[8] & B[1]), .ci(carry1[7]), .s(sum1[8]), .co(carry1[8]));
FA fa1_9(.a(sum0[10]), .b(A[9] & B[1]), .ci(carry1[8]), .s(sum1[9]), .co(carry1[9]));
FA fa1_10(.a(sum0[11]), .b(A[10] & B[1]), .ci(carry1[9]), .s(sum1[10]), .co(carry1[10]));
FA fa1_11(.a(sum0[12]), .b(A[11] & B[1]), .ci(carry1[10]), .s(sum1[11]), .co(carry1[11]));
FA fa1_12(.a(sum0[13]), .b(A[12] & B[1]), .ci(carry1[11]), .s(sum1[12]), .co(carry1[12]));
FA fa1_13(.a(sum0[14]), .b(A[13] & B[1]), .ci(carry1[12]), .s(sum1[13]), .co(carry1[13]));
FA fa1_14(.a(sum0[15]), .b(A[14] & B[1]), .ci(carry1[13]), .s(sum1[14]), .co(carry1[14]));
FA fa1_15(.a(sum0[16]), .b(A[15] & B[1]), .ci(carry1[14]), .s(sum1[15]), .co(carry1[15]));
FA fa1_16(.a(sum0[17]), .b(A[16] & B[1]), .ci(carry1[15]), .s(sum1[16]), .co(carry1[16]));
FA fa1_17(.a(sum0[18]), .b(A[17] & B[1]), .ci(carry1[16]), .s(sum1[17]), .co(carry1[17]));
FA fa1_18(.a(sum0[19]), .b(A[18] & B[1]), .ci(carry1[17]), .s(sum1[18]), .co(carry1[18]));
FA fa1_19(.a(sum0[20]), .b(A[19] & B[1]), .ci(carry1[18]), .s(sum1[19]), .co(carry1[19]));
FA fa1_20(.a(sum0[21]), .b(A[20] & B[1]), .ci(carry1[19]), .s(sum1[20]), .co(carry1[20]));
FA fa1_21(.a(sum0[22]), .b(A[21] & B[1]), .ci(carry1[20]), .s(sum1[21]), .co(carry1[21]));
FA fa1_22(.a(sum0[23]), .b(A[22] & B[1]), .ci(carry1[21]), .s(sum1[22]), .co(carry1[22]));
FA fa1_23(.a(sum0[24]), .b(A[23] & B[1]), .ci(carry1[22]), .s(sum1[23]), .co(carry1[23]));
FA fa1_24(.a(sum0[25]), .b(A[24] & B[1]), .ci(carry1[23]), .s(sum1[24]), .co(carry1[24]));
FA fa1_25(.a(sum0[26]), .b(A[25] & B[1]), .ci(carry1[24]), .s(sum1[25]), .co(carry1[25]));
FA fa1_26(.a(sum0[27]), .b(A[26] & B[1]), .ci(carry1[25]), .s(sum1[26]), .co(carry1[26]));
FA fa1_27(.a(sum0[28]), .b(A[27] & B[1]), .ci(carry1[26]), .s(sum1[27]), .co(carry1[27]));
FA fa1_28(.a(sum0[29]), .b(A[28] & B[1]), .ci(carry1[27]), .s(sum1[28]), .co(carry1[28]));
FA fa1_29(.a(sum0[30]), .b(A[29] & B[1]), .ci(carry1[28]), .s(sum1[29]), .co(carry1[29]));
FA fa1_30(.a(sum0[31]), .b(A[30] & B[1]), .ci(carry1[29]), .s(sum1[30]), .co(carry1[30]));
FA fa1_31(.a(carry0[31]), .b(A[31] & B[1]), .ci(carry1[30]), .s(sum1[31]), .co(carry1[31]));
FA fa2_0(.a(sum1[1]), .b(A[0] & B[2]), .ci(1'b0), .s(Z[2]), .co(carry2[0]));
FA fa2_1(.a(sum1[2]), .b(A[1] & B[2]), .ci(carry2[0]), .s(sum2[1]), .co(carry2[1]));
FA fa2_2(.a(sum1[3]), .b(A[2] & B[2]), .ci(carry2[1]), .s(sum2[2]), .co(carry2[2]));
FA fa2_3(.a(sum1[4]), .b(A[3] & B[2]), .ci(carry2[2]), .s(sum2[3]), .co(carry2[3]));
FA fa2_4(.a(sum1[5]), .b(A[4] & B[2]), .ci(carry2[3]), .s(sum2[4]), .co(carry2[4]));
FA fa2_5(.a(sum1[6]), .b(A[5] & B[2]), .ci(carry2[4]), .s(sum2[5]), .co(carry2[5]));
FA fa2_6(.a(sum1[7]), .b(A[6] & B[2]), .ci(carry2[5]), .s(sum2[6]), .co(carry2[6]));
FA fa2_7(.a(sum1[8]), .b(A[7] & B[2]), .ci(carry2[6]), .s(sum2[7]), .co(carry2[7]));
FA fa2_8(.a(sum1[9]), .b(A[8] & B[2]), .ci(carry2[7]), .s(sum2[8]), .co(carry2[8]));
FA fa2_9(.a(sum1[10]), .b(A[9] & B[2]), .ci(carry2[8]), .s(sum2[9]), .co(carry2[9]));
FA fa2_10(.a(sum1[11]), .b(A[10] & B[2]), .ci(carry2[9]), .s(sum2[10]), .co(carry2[10]));
FA fa2_11(.a(sum1[12]), .b(A[11] & B[2]), .ci(carry2[10]), .s(sum2[11]), .co(carry2[11]));
FA fa2_12(.a(sum1[13]), .b(A[12] & B[2]), .ci(carry2[11]), .s(sum2[12]), .co(carry2[12]));
FA fa2_13(.a(sum1[14]), .b(A[13] & B[2]), .ci(carry2[12]), .s(sum2[13]), .co(carry2[13]));
FA fa2_14(.a(sum1[15]), .b(A[14] & B[2]), .ci(carry2[13]), .s(sum2[14]), .co(carry2[14]));
FA fa2_15(.a(sum1[16]), .b(A[15] & B[2]), .ci(carry2[14]), .s(sum2[15]), .co(carry2[15]));
FA fa2_16(.a(sum1[17]), .b(A[16] & B[2]), .ci(carry2[15]), .s(sum2[16]), .co(carry2[16]));
FA fa2_17(.a(sum1[18]), .b(A[17] & B[2]), .ci(carry2[16]), .s(sum2[17]), .co(carry2[17]));
FA fa2_18(.a(sum1[19]), .b(A[18] & B[2]), .ci(carry2[17]), .s(sum2[18]), .co(carry2[18]));
FA fa2_19(.a(sum1[20]), .b(A[19] & B[2]), .ci(carry2[18]), .s(sum2[19]), .co(carry2[19]));
FA fa2_20(.a(sum1[21]), .b(A[20] & B[2]), .ci(carry2[19]), .s(sum2[20]), .co(carry2[20]));
FA fa2_21(.a(sum1[22]), .b(A[21] & B[2]), .ci(carry2[20]), .s(sum2[21]), .co(carry2[21]));
FA fa2_22(.a(sum1[23]), .b(A[22] & B[2]), .ci(carry2[21]), .s(sum2[22]), .co(carry2[22]));
FA fa2_23(.a(sum1[24]), .b(A[23] & B[2]), .ci(carry2[22]), .s(sum2[23]), .co(carry2[23]));
FA fa2_24(.a(sum1[25]), .b(A[24] & B[2]), .ci(carry2[23]), .s(sum2[24]), .co(carry2[24]));
FA fa2_25(.a(sum1[26]), .b(A[25] & B[2]), .ci(carry2[24]), .s(sum2[25]), .co(carry2[25]));
FA fa2_26(.a(sum1[27]), .b(A[26] & B[2]), .ci(carry2[25]), .s(sum2[26]), .co(carry2[26]));
FA fa2_27(.a(sum1[28]), .b(A[27] & B[2]), .ci(carry2[26]), .s(sum2[27]), .co(carry2[27]));
FA fa2_28(.a(sum1[29]), .b(A[28] & B[2]), .ci(carry2[27]), .s(sum2[28]), .co(carry2[28]));
FA fa2_29(.a(sum1[30]), .b(A[29] & B[2]), .ci(carry2[28]), .s(sum2[29]), .co(carry2[29]));
FA fa2_30(.a(sum1[31]), .b(A[30] & B[2]), .ci(carry2[29]), .s(sum2[30]), .co(carry2[30]));
FA fa2_31(.a(carry1[31]), .b(A[31] & B[2]), .ci(carry2[30]), .s(sum2[31]), .co(carry2[31]));
FA fa3_0(.a(sum2[1]), .b(A[0] & B[3]), .ci(1'b0), .s(Z[3]), .co(carry3[0]));
FA fa3_1(.a(sum2[2]), .b(A[1] & B[3]), .ci(carry3[0]), .s(sum3[1]), .co(carry3[1]));
FA fa3_2(.a(sum2[3]), .b(A[2] & B[3]), .ci(carry3[1]), .s(sum3[2]), .co(carry3[2]));
FA fa3_3(.a(sum2[4]), .b(A[3] & B[3]), .ci(carry3[2]), .s(sum3[3]), .co(carry3[3]));
FA fa3_4(.a(sum2[5]), .b(A[4] & B[3]), .ci(carry3[3]), .s(sum3[4]), .co(carry3[4]));
FA fa3_5(.a(sum2[6]), .b(A[5] & B[3]), .ci(carry3[4]), .s(sum3[5]), .co(carry3[5]));
FA fa3_6(.a(sum2[7]), .b(A[6] & B[3]), .ci(carry3[5]), .s(sum3[6]), .co(carry3[6]));
FA fa3_7(.a(sum2[8]), .b(A[7] & B[3]), .ci(carry3[6]), .s(sum3[7]), .co(carry3[7]));
FA fa3_8(.a(sum2[9]), .b(A[8] & B[3]), .ci(carry3[7]), .s(sum3[8]), .co(carry3[8]));
FA fa3_9(.a(sum2[10]), .b(A[9] & B[3]), .ci(carry3[8]), .s(sum3[9]), .co(carry3[9]));
FA fa3_10(.a(sum2[11]), .b(A[10] & B[3]), .ci(carry3[9]), .s(sum3[10]), .co(carry3[10]));
FA fa3_11(.a(sum2[12]), .b(A[11] & B[3]), .ci(carry3[10]), .s(sum3[11]), .co(carry3[11]));
FA fa3_12(.a(sum2[13]), .b(A[12] & B[3]), .ci(carry3[11]), .s(sum3[12]), .co(carry3[12]));
FA fa3_13(.a(sum2[14]), .b(A[13] & B[3]), .ci(carry3[12]), .s(sum3[13]), .co(carry3[13]));
FA fa3_14(.a(sum2[15]), .b(A[14] & B[3]), .ci(carry3[13]), .s(sum3[14]), .co(carry3[14]));
FA fa3_15(.a(sum2[16]), .b(A[15] & B[3]), .ci(carry3[14]), .s(sum3[15]), .co(carry3[15]));
FA fa3_16(.a(sum2[17]), .b(A[16] & B[3]), .ci(carry3[15]), .s(sum3[16]), .co(carry3[16]));
FA fa3_17(.a(sum2[18]), .b(A[17] & B[3]), .ci(carry3[16]), .s(sum3[17]), .co(carry3[17]));
FA fa3_18(.a(sum2[19]), .b(A[18] & B[3]), .ci(carry3[17]), .s(sum3[18]), .co(carry3[18]));
FA fa3_19(.a(sum2[20]), .b(A[19] & B[3]), .ci(carry3[18]), .s(sum3[19]), .co(carry3[19]));
FA fa3_20(.a(sum2[21]), .b(A[20] & B[3]), .ci(carry3[19]), .s(sum3[20]), .co(carry3[20]));
FA fa3_21(.a(sum2[22]), .b(A[21] & B[3]), .ci(carry3[20]), .s(sum3[21]), .co(carry3[21]));
FA fa3_22(.a(sum2[23]), .b(A[22] & B[3]), .ci(carry3[21]), .s(sum3[22]), .co(carry3[22]));
FA fa3_23(.a(sum2[24]), .b(A[23] & B[3]), .ci(carry3[22]), .s(sum3[23]), .co(carry3[23]));
FA fa3_24(.a(sum2[25]), .b(A[24] & B[3]), .ci(carry3[23]), .s(sum3[24]), .co(carry3[24]));
FA fa3_25(.a(sum2[26]), .b(A[25] & B[3]), .ci(carry3[24]), .s(sum3[25]), .co(carry3[25]));
FA fa3_26(.a(sum2[27]), .b(A[26] & B[3]), .ci(carry3[25]), .s(sum3[26]), .co(carry3[26]));
FA fa3_27(.a(sum2[28]), .b(A[27] & B[3]), .ci(carry3[26]), .s(sum3[27]), .co(carry3[27]));
FA fa3_28(.a(sum2[29]), .b(A[28] & B[3]), .ci(carry3[27]), .s(sum3[28]), .co(carry3[28]));
FA fa3_29(.a(sum2[30]), .b(A[29] & B[3]), .ci(carry3[28]), .s(sum3[29]), .co(carry3[29]));
FA fa3_30(.a(sum2[31]), .b(A[30] & B[3]), .ci(carry3[29]), .s(sum3[30]), .co(carry3[30]));
FA fa3_31(.a(carry2[31]), .b(A[31] & B[3]), .ci(carry3[30]), .s(sum3[31]), .co(carry3[31]));
FA fa4_0(.a(sum3[1]), .b(A[0] & B[4]), .ci(1'b0), .s(Z[4]), .co(carry4[0]));
FA fa4_1(.a(sum3[2]), .b(A[1] & B[4]), .ci(carry4[0]), .s(sum4[1]), .co(carry4[1]));
FA fa4_2(.a(sum3[3]), .b(A[2] & B[4]), .ci(carry4[1]), .s(sum4[2]), .co(carry4[2]));
FA fa4_3(.a(sum3[4]), .b(A[3] & B[4]), .ci(carry4[2]), .s(sum4[3]), .co(carry4[3]));
FA fa4_4(.a(sum3[5]), .b(A[4] & B[4]), .ci(carry4[3]), .s(sum4[4]), .co(carry4[4]));
FA fa4_5(.a(sum3[6]), .b(A[5] & B[4]), .ci(carry4[4]), .s(sum4[5]), .co(carry4[5]));
FA fa4_6(.a(sum3[7]), .b(A[6] & B[4]), .ci(carry4[5]), .s(sum4[6]), .co(carry4[6]));
FA fa4_7(.a(sum3[8]), .b(A[7] & B[4]), .ci(carry4[6]), .s(sum4[7]), .co(carry4[7]));
FA fa4_8(.a(sum3[9]), .b(A[8] & B[4]), .ci(carry4[7]), .s(sum4[8]), .co(carry4[8]));
FA fa4_9(.a(sum3[10]), .b(A[9] & B[4]), .ci(carry4[8]), .s(sum4[9]), .co(carry4[9]));
FA fa4_10(.a(sum3[11]), .b(A[10] & B[4]), .ci(carry4[9]), .s(sum4[10]), .co(carry4[10]));
FA fa4_11(.a(sum3[12]), .b(A[11] & B[4]), .ci(carry4[10]), .s(sum4[11]), .co(carry4[11]));
FA fa4_12(.a(sum3[13]), .b(A[12] & B[4]), .ci(carry4[11]), .s(sum4[12]), .co(carry4[12]));
FA fa4_13(.a(sum3[14]), .b(A[13] & B[4]), .ci(carry4[12]), .s(sum4[13]), .co(carry4[13]));
FA fa4_14(.a(sum3[15]), .b(A[14] & B[4]), .ci(carry4[13]), .s(sum4[14]), .co(carry4[14]));
FA fa4_15(.a(sum3[16]), .b(A[15] & B[4]), .ci(carry4[14]), .s(sum4[15]), .co(carry4[15]));
FA fa4_16(.a(sum3[17]), .b(A[16] & B[4]), .ci(carry4[15]), .s(sum4[16]), .co(carry4[16]));
FA fa4_17(.a(sum3[18]), .b(A[17] & B[4]), .ci(carry4[16]), .s(sum4[17]), .co(carry4[17]));
FA fa4_18(.a(sum3[19]), .b(A[18] & B[4]), .ci(carry4[17]), .s(sum4[18]), .co(carry4[18]));
FA fa4_19(.a(sum3[20]), .b(A[19] & B[4]), .ci(carry4[18]), .s(sum4[19]), .co(carry4[19]));
FA fa4_20(.a(sum3[21]), .b(A[20] & B[4]), .ci(carry4[19]), .s(sum4[20]), .co(carry4[20]));
FA fa4_21(.a(sum3[22]), .b(A[21] & B[4]), .ci(carry4[20]), .s(sum4[21]), .co(carry4[21]));
FA fa4_22(.a(sum3[23]), .b(A[22] & B[4]), .ci(carry4[21]), .s(sum4[22]), .co(carry4[22]));
FA fa4_23(.a(sum3[24]), .b(A[23] & B[4]), .ci(carry4[22]), .s(sum4[23]), .co(carry4[23]));
FA fa4_24(.a(sum3[25]), .b(A[24] & B[4]), .ci(carry4[23]), .s(sum4[24]), .co(carry4[24]));
FA fa4_25(.a(sum3[26]), .b(A[25] & B[4]), .ci(carry4[24]), .s(sum4[25]), .co(carry4[25]));
FA fa4_26(.a(sum3[27]), .b(A[26] & B[4]), .ci(carry4[25]), .s(sum4[26]), .co(carry4[26]));
FA fa4_27(.a(sum3[28]), .b(A[27] & B[4]), .ci(carry4[26]), .s(sum4[27]), .co(carry4[27]));
FA fa4_28(.a(sum3[29]), .b(A[28] & B[4]), .ci(carry4[27]), .s(sum4[28]), .co(carry4[28]));
FA fa4_29(.a(sum3[30]), .b(A[29] & B[4]), .ci(carry4[28]), .s(sum4[29]), .co(carry4[29]));
FA fa4_30(.a(sum3[31]), .b(A[30] & B[4]), .ci(carry4[29]), .s(sum4[30]), .co(carry4[30]));
FA fa4_31(.a(carry3[31]), .b(A[31] & B[4]), .ci(carry4[30]), .s(sum4[31]), .co(carry4[31]));
FA fa5_0(.a(sum4[1]), .b(A[0] & B[5]), .ci(1'b0), .s(Z[5]), .co(carry5[0]));
FA fa5_1(.a(sum4[2]), .b(A[1] & B[5]), .ci(carry5[0]), .s(sum5[1]), .co(carry5[1]));
FA fa5_2(.a(sum4[3]), .b(A[2] & B[5]), .ci(carry5[1]), .s(sum5[2]), .co(carry5[2]));
FA fa5_3(.a(sum4[4]), .b(A[3] & B[5]), .ci(carry5[2]), .s(sum5[3]), .co(carry5[3]));
FA fa5_4(.a(sum4[5]), .b(A[4] & B[5]), .ci(carry5[3]), .s(sum5[4]), .co(carry5[4]));
FA fa5_5(.a(sum4[6]), .b(A[5] & B[5]), .ci(carry5[4]), .s(sum5[5]), .co(carry5[5]));
FA fa5_6(.a(sum4[7]), .b(A[6] & B[5]), .ci(carry5[5]), .s(sum5[6]), .co(carry5[6]));
FA fa5_7(.a(sum4[8]), .b(A[7] & B[5]), .ci(carry5[6]), .s(sum5[7]), .co(carry5[7]));
FA fa5_8(.a(sum4[9]), .b(A[8] & B[5]), .ci(carry5[7]), .s(sum5[8]), .co(carry5[8]));
FA fa5_9(.a(sum4[10]), .b(A[9] & B[5]), .ci(carry5[8]), .s(sum5[9]), .co(carry5[9]));
FA fa5_10(.a(sum4[11]), .b(A[10] & B[5]), .ci(carry5[9]), .s(sum5[10]), .co(carry5[10]));
FA fa5_11(.a(sum4[12]), .b(A[11] & B[5]), .ci(carry5[10]), .s(sum5[11]), .co(carry5[11]));
FA fa5_12(.a(sum4[13]), .b(A[12] & B[5]), .ci(carry5[11]), .s(sum5[12]), .co(carry5[12]));
FA fa5_13(.a(sum4[14]), .b(A[13] & B[5]), .ci(carry5[12]), .s(sum5[13]), .co(carry5[13]));
FA fa5_14(.a(sum4[15]), .b(A[14] & B[5]), .ci(carry5[13]), .s(sum5[14]), .co(carry5[14]));
FA fa5_15(.a(sum4[16]), .b(A[15] & B[5]), .ci(carry5[14]), .s(sum5[15]), .co(carry5[15]));
FA fa5_16(.a(sum4[17]), .b(A[16] & B[5]), .ci(carry5[15]), .s(sum5[16]), .co(carry5[16]));
FA fa5_17(.a(sum4[18]), .b(A[17] & B[5]), .ci(carry5[16]), .s(sum5[17]), .co(carry5[17]));
FA fa5_18(.a(sum4[19]), .b(A[18] & B[5]), .ci(carry5[17]), .s(sum5[18]), .co(carry5[18]));
FA fa5_19(.a(sum4[20]), .b(A[19] & B[5]), .ci(carry5[18]), .s(sum5[19]), .co(carry5[19]));
FA fa5_20(.a(sum4[21]), .b(A[20] & B[5]), .ci(carry5[19]), .s(sum5[20]), .co(carry5[20]));
FA fa5_21(.a(sum4[22]), .b(A[21] & B[5]), .ci(carry5[20]), .s(sum5[21]), .co(carry5[21]));
FA fa5_22(.a(sum4[23]), .b(A[22] & B[5]), .ci(carry5[21]), .s(sum5[22]), .co(carry5[22]));
FA fa5_23(.a(sum4[24]), .b(A[23] & B[5]), .ci(carry5[22]), .s(sum5[23]), .co(carry5[23]));
FA fa5_24(.a(sum4[25]), .b(A[24] & B[5]), .ci(carry5[23]), .s(sum5[24]), .co(carry5[24]));
FA fa5_25(.a(sum4[26]), .b(A[25] & B[5]), .ci(carry5[24]), .s(sum5[25]), .co(carry5[25]));
FA fa5_26(.a(sum4[27]), .b(A[26] & B[5]), .ci(carry5[25]), .s(sum5[26]), .co(carry5[26]));
FA fa5_27(.a(sum4[28]), .b(A[27] & B[5]), .ci(carry5[26]), .s(sum5[27]), .co(carry5[27]));
FA fa5_28(.a(sum4[29]), .b(A[28] & B[5]), .ci(carry5[27]), .s(sum5[28]), .co(carry5[28]));
FA fa5_29(.a(sum4[30]), .b(A[29] & B[5]), .ci(carry5[28]), .s(sum5[29]), .co(carry5[29]));
FA fa5_30(.a(sum4[31]), .b(A[30] & B[5]), .ci(carry5[29]), .s(sum5[30]), .co(carry5[30]));
FA fa5_31(.a(carry4[31]), .b(A[31] & B[5]), .ci(carry5[30]), .s(sum5[31]), .co(carry5[31]));
FA fa6_0(.a(sum5[1]), .b(A[0] & B[6]), .ci(1'b0), .s(Z[6]), .co(carry6[0]));
FA fa6_1(.a(sum5[2]), .b(A[1] & B[6]), .ci(carry6[0]), .s(sum6[1]), .co(carry6[1]));
FA fa6_2(.a(sum5[3]), .b(A[2] & B[6]), .ci(carry6[1]), .s(sum6[2]), .co(carry6[2]));
FA fa6_3(.a(sum5[4]), .b(A[3] & B[6]), .ci(carry6[2]), .s(sum6[3]), .co(carry6[3]));
FA fa6_4(.a(sum5[5]), .b(A[4] & B[6]), .ci(carry6[3]), .s(sum6[4]), .co(carry6[4]));
FA fa6_5(.a(sum5[6]), .b(A[5] & B[6]), .ci(carry6[4]), .s(sum6[5]), .co(carry6[5]));
FA fa6_6(.a(sum5[7]), .b(A[6] & B[6]), .ci(carry6[5]), .s(sum6[6]), .co(carry6[6]));
FA fa6_7(.a(sum5[8]), .b(A[7] & B[6]), .ci(carry6[6]), .s(sum6[7]), .co(carry6[7]));
FA fa6_8(.a(sum5[9]), .b(A[8] & B[6]), .ci(carry6[7]), .s(sum6[8]), .co(carry6[8]));
FA fa6_9(.a(sum5[10]), .b(A[9] & B[6]), .ci(carry6[8]), .s(sum6[9]), .co(carry6[9]));
FA fa6_10(.a(sum5[11]), .b(A[10] & B[6]), .ci(carry6[9]), .s(sum6[10]), .co(carry6[10]));
FA fa6_11(.a(sum5[12]), .b(A[11] & B[6]), .ci(carry6[10]), .s(sum6[11]), .co(carry6[11]));
FA fa6_12(.a(sum5[13]), .b(A[12] & B[6]), .ci(carry6[11]), .s(sum6[12]), .co(carry6[12]));
FA fa6_13(.a(sum5[14]), .b(A[13] & B[6]), .ci(carry6[12]), .s(sum6[13]), .co(carry6[13]));
FA fa6_14(.a(sum5[15]), .b(A[14] & B[6]), .ci(carry6[13]), .s(sum6[14]), .co(carry6[14]));
FA fa6_15(.a(sum5[16]), .b(A[15] & B[6]), .ci(carry6[14]), .s(sum6[15]), .co(carry6[15]));
FA fa6_16(.a(sum5[17]), .b(A[16] & B[6]), .ci(carry6[15]), .s(sum6[16]), .co(carry6[16]));
FA fa6_17(.a(sum5[18]), .b(A[17] & B[6]), .ci(carry6[16]), .s(sum6[17]), .co(carry6[17]));
FA fa6_18(.a(sum5[19]), .b(A[18] & B[6]), .ci(carry6[17]), .s(sum6[18]), .co(carry6[18]));
FA fa6_19(.a(sum5[20]), .b(A[19] & B[6]), .ci(carry6[18]), .s(sum6[19]), .co(carry6[19]));
FA fa6_20(.a(sum5[21]), .b(A[20] & B[6]), .ci(carry6[19]), .s(sum6[20]), .co(carry6[20]));
FA fa6_21(.a(sum5[22]), .b(A[21] & B[6]), .ci(carry6[20]), .s(sum6[21]), .co(carry6[21]));
FA fa6_22(.a(sum5[23]), .b(A[22] & B[6]), .ci(carry6[21]), .s(sum6[22]), .co(carry6[22]));
FA fa6_23(.a(sum5[24]), .b(A[23] & B[6]), .ci(carry6[22]), .s(sum6[23]), .co(carry6[23]));
FA fa6_24(.a(sum5[25]), .b(A[24] & B[6]), .ci(carry6[23]), .s(sum6[24]), .co(carry6[24]));
FA fa6_25(.a(sum5[26]), .b(A[25] & B[6]), .ci(carry6[24]), .s(sum6[25]), .co(carry6[25]));
FA fa6_26(.a(sum5[27]), .b(A[26] & B[6]), .ci(carry6[25]), .s(sum6[26]), .co(carry6[26]));
FA fa6_27(.a(sum5[28]), .b(A[27] & B[6]), .ci(carry6[26]), .s(sum6[27]), .co(carry6[27]));
FA fa6_28(.a(sum5[29]), .b(A[28] & B[6]), .ci(carry6[27]), .s(sum6[28]), .co(carry6[28]));
FA fa6_29(.a(sum5[30]), .b(A[29] & B[6]), .ci(carry6[28]), .s(sum6[29]), .co(carry6[29]));
FA fa6_30(.a(sum5[31]), .b(A[30] & B[6]), .ci(carry6[29]), .s(sum6[30]), .co(carry6[30]));
FA fa6_31(.a(carry5[31]), .b(A[31] & B[6]), .ci(carry6[30]), .s(sum6[31]), .co(carry6[31]));
FA fa7_0(.a(sum6[1]), .b(A[0] & B[7]), .ci(1'b0), .s(Z[7]), .co(carry7[0]));
FA fa7_1(.a(sum6[2]), .b(A[1] & B[7]), .ci(carry7[0]), .s(sum7[1]), .co(carry7[1]));
FA fa7_2(.a(sum6[3]), .b(A[2] & B[7]), .ci(carry7[1]), .s(sum7[2]), .co(carry7[2]));
FA fa7_3(.a(sum6[4]), .b(A[3] & B[7]), .ci(carry7[2]), .s(sum7[3]), .co(carry7[3]));
FA fa7_4(.a(sum6[5]), .b(A[4] & B[7]), .ci(carry7[3]), .s(sum7[4]), .co(carry7[4]));
FA fa7_5(.a(sum6[6]), .b(A[5] & B[7]), .ci(carry7[4]), .s(sum7[5]), .co(carry7[5]));
FA fa7_6(.a(sum6[7]), .b(A[6] & B[7]), .ci(carry7[5]), .s(sum7[6]), .co(carry7[6]));
FA fa7_7(.a(sum6[8]), .b(A[7] & B[7]), .ci(carry7[6]), .s(sum7[7]), .co(carry7[7]));
FA fa7_8(.a(sum6[9]), .b(A[8] & B[7]), .ci(carry7[7]), .s(sum7[8]), .co(carry7[8]));
FA fa7_9(.a(sum6[10]), .b(A[9] & B[7]), .ci(carry7[8]), .s(sum7[9]), .co(carry7[9]));
FA fa7_10(.a(sum6[11]), .b(A[10] & B[7]), .ci(carry7[9]), .s(sum7[10]), .co(carry7[10]));
FA fa7_11(.a(sum6[12]), .b(A[11] & B[7]), .ci(carry7[10]), .s(sum7[11]), .co(carry7[11]));
FA fa7_12(.a(sum6[13]), .b(A[12] & B[7]), .ci(carry7[11]), .s(sum7[12]), .co(carry7[12]));
FA fa7_13(.a(sum6[14]), .b(A[13] & B[7]), .ci(carry7[12]), .s(sum7[13]), .co(carry7[13]));
FA fa7_14(.a(sum6[15]), .b(A[14] & B[7]), .ci(carry7[13]), .s(sum7[14]), .co(carry7[14]));
FA fa7_15(.a(sum6[16]), .b(A[15] & B[7]), .ci(carry7[14]), .s(sum7[15]), .co(carry7[15]));
FA fa7_16(.a(sum6[17]), .b(A[16] & B[7]), .ci(carry7[15]), .s(sum7[16]), .co(carry7[16]));
FA fa7_17(.a(sum6[18]), .b(A[17] & B[7]), .ci(carry7[16]), .s(sum7[17]), .co(carry7[17]));
FA fa7_18(.a(sum6[19]), .b(A[18] & B[7]), .ci(carry7[17]), .s(sum7[18]), .co(carry7[18]));
FA fa7_19(.a(sum6[20]), .b(A[19] & B[7]), .ci(carry7[18]), .s(sum7[19]), .co(carry7[19]));
FA fa7_20(.a(sum6[21]), .b(A[20] & B[7]), .ci(carry7[19]), .s(sum7[20]), .co(carry7[20]));
FA fa7_21(.a(sum6[22]), .b(A[21] & B[7]), .ci(carry7[20]), .s(sum7[21]), .co(carry7[21]));
FA fa7_22(.a(sum6[23]), .b(A[22] & B[7]), .ci(carry7[21]), .s(sum7[22]), .co(carry7[22]));
FA fa7_23(.a(sum6[24]), .b(A[23] & B[7]), .ci(carry7[22]), .s(sum7[23]), .co(carry7[23]));
FA fa7_24(.a(sum6[25]), .b(A[24] & B[7]), .ci(carry7[23]), .s(sum7[24]), .co(carry7[24]));
FA fa7_25(.a(sum6[26]), .b(A[25] & B[7]), .ci(carry7[24]), .s(sum7[25]), .co(carry7[25]));
FA fa7_26(.a(sum6[27]), .b(A[26] & B[7]), .ci(carry7[25]), .s(sum7[26]), .co(carry7[26]));
FA fa7_27(.a(sum6[28]), .b(A[27] & B[7]), .ci(carry7[26]), .s(sum7[27]), .co(carry7[27]));
FA fa7_28(.a(sum6[29]), .b(A[28] & B[7]), .ci(carry7[27]), .s(sum7[28]), .co(carry7[28]));
FA fa7_29(.a(sum6[30]), .b(A[29] & B[7]), .ci(carry7[28]), .s(sum7[29]), .co(carry7[29]));
FA fa7_30(.a(sum6[31]), .b(A[30] & B[7]), .ci(carry7[29]), .s(sum7[30]), .co(carry7[30]));
FA fa7_31(.a(carry6[31]), .b(A[31] & B[7]), .ci(carry7[30]), .s(sum7[31]), .co(carry7[31]));
FA fa8_0(.a(sum7[1]), .b(A[0] & B[8]), .ci(1'b0), .s(Z[8]), .co(carry8[0]));
FA fa8_1(.a(sum7[2]), .b(A[1] & B[8]), .ci(carry8[0]), .s(sum8[1]), .co(carry8[1]));
FA fa8_2(.a(sum7[3]), .b(A[2] & B[8]), .ci(carry8[1]), .s(sum8[2]), .co(carry8[2]));
FA fa8_3(.a(sum7[4]), .b(A[3] & B[8]), .ci(carry8[2]), .s(sum8[3]), .co(carry8[3]));
FA fa8_4(.a(sum7[5]), .b(A[4] & B[8]), .ci(carry8[3]), .s(sum8[4]), .co(carry8[4]));
FA fa8_5(.a(sum7[6]), .b(A[5] & B[8]), .ci(carry8[4]), .s(sum8[5]), .co(carry8[5]));
FA fa8_6(.a(sum7[7]), .b(A[6] & B[8]), .ci(carry8[5]), .s(sum8[6]), .co(carry8[6]));
FA fa8_7(.a(sum7[8]), .b(A[7] & B[8]), .ci(carry8[6]), .s(sum8[7]), .co(carry8[7]));
FA fa8_8(.a(sum7[9]), .b(A[8] & B[8]), .ci(carry8[7]), .s(sum8[8]), .co(carry8[8]));
FA fa8_9(.a(sum7[10]), .b(A[9] & B[8]), .ci(carry8[8]), .s(sum8[9]), .co(carry8[9]));
FA fa8_10(.a(sum7[11]), .b(A[10] & B[8]), .ci(carry8[9]), .s(sum8[10]), .co(carry8[10]));
FA fa8_11(.a(sum7[12]), .b(A[11] & B[8]), .ci(carry8[10]), .s(sum8[11]), .co(carry8[11]));
FA fa8_12(.a(sum7[13]), .b(A[12] & B[8]), .ci(carry8[11]), .s(sum8[12]), .co(carry8[12]));
FA fa8_13(.a(sum7[14]), .b(A[13] & B[8]), .ci(carry8[12]), .s(sum8[13]), .co(carry8[13]));
FA fa8_14(.a(sum7[15]), .b(A[14] & B[8]), .ci(carry8[13]), .s(sum8[14]), .co(carry8[14]));
FA fa8_15(.a(sum7[16]), .b(A[15] & B[8]), .ci(carry8[14]), .s(sum8[15]), .co(carry8[15]));
FA fa8_16(.a(sum7[17]), .b(A[16] & B[8]), .ci(carry8[15]), .s(sum8[16]), .co(carry8[16]));
FA fa8_17(.a(sum7[18]), .b(A[17] & B[8]), .ci(carry8[16]), .s(sum8[17]), .co(carry8[17]));
FA fa8_18(.a(sum7[19]), .b(A[18] & B[8]), .ci(carry8[17]), .s(sum8[18]), .co(carry8[18]));
FA fa8_19(.a(sum7[20]), .b(A[19] & B[8]), .ci(carry8[18]), .s(sum8[19]), .co(carry8[19]));
FA fa8_20(.a(sum7[21]), .b(A[20] & B[8]), .ci(carry8[19]), .s(sum8[20]), .co(carry8[20]));
FA fa8_21(.a(sum7[22]), .b(A[21] & B[8]), .ci(carry8[20]), .s(sum8[21]), .co(carry8[21]));
FA fa8_22(.a(sum7[23]), .b(A[22] & B[8]), .ci(carry8[21]), .s(sum8[22]), .co(carry8[22]));
FA fa8_23(.a(sum7[24]), .b(A[23] & B[8]), .ci(carry8[22]), .s(sum8[23]), .co(carry8[23]));
FA fa8_24(.a(sum7[25]), .b(A[24] & B[8]), .ci(carry8[23]), .s(sum8[24]), .co(carry8[24]));
FA fa8_25(.a(sum7[26]), .b(A[25] & B[8]), .ci(carry8[24]), .s(sum8[25]), .co(carry8[25]));
FA fa8_26(.a(sum7[27]), .b(A[26] & B[8]), .ci(carry8[25]), .s(sum8[26]), .co(carry8[26]));
FA fa8_27(.a(sum7[28]), .b(A[27] & B[8]), .ci(carry8[26]), .s(sum8[27]), .co(carry8[27]));
FA fa8_28(.a(sum7[29]), .b(A[28] & B[8]), .ci(carry8[27]), .s(sum8[28]), .co(carry8[28]));
FA fa8_29(.a(sum7[30]), .b(A[29] & B[8]), .ci(carry8[28]), .s(sum8[29]), .co(carry8[29]));
FA fa8_30(.a(sum7[31]), .b(A[30] & B[8]), .ci(carry8[29]), .s(sum8[30]), .co(carry8[30]));
FA fa8_31(.a(carry7[31]), .b(A[31] & B[8]), .ci(carry8[30]), .s(sum8[31]), .co(carry8[31]));
FA fa9_0(.a(sum8[1]), .b(A[0] & B[9]), .ci(1'b0), .s(Z[9]), .co(carry9[0]));
FA fa9_1(.a(sum8[2]), .b(A[1] & B[9]), .ci(carry9[0]), .s(sum9[1]), .co(carry9[1]));
FA fa9_2(.a(sum8[3]), .b(A[2] & B[9]), .ci(carry9[1]), .s(sum9[2]), .co(carry9[2]));
FA fa9_3(.a(sum8[4]), .b(A[3] & B[9]), .ci(carry9[2]), .s(sum9[3]), .co(carry9[3]));
FA fa9_4(.a(sum8[5]), .b(A[4] & B[9]), .ci(carry9[3]), .s(sum9[4]), .co(carry9[4]));
FA fa9_5(.a(sum8[6]), .b(A[5] & B[9]), .ci(carry9[4]), .s(sum9[5]), .co(carry9[5]));
FA fa9_6(.a(sum8[7]), .b(A[6] & B[9]), .ci(carry9[5]), .s(sum9[6]), .co(carry9[6]));
FA fa9_7(.a(sum8[8]), .b(A[7] & B[9]), .ci(carry9[6]), .s(sum9[7]), .co(carry9[7]));
FA fa9_8(.a(sum8[9]), .b(A[8] & B[9]), .ci(carry9[7]), .s(sum9[8]), .co(carry9[8]));
FA fa9_9(.a(sum8[10]), .b(A[9] & B[9]), .ci(carry9[8]), .s(sum9[9]), .co(carry9[9]));
FA fa9_10(.a(sum8[11]), .b(A[10] & B[9]), .ci(carry9[9]), .s(sum9[10]), .co(carry9[10]));
FA fa9_11(.a(sum8[12]), .b(A[11] & B[9]), .ci(carry9[10]), .s(sum9[11]), .co(carry9[11]));
FA fa9_12(.a(sum8[13]), .b(A[12] & B[9]), .ci(carry9[11]), .s(sum9[12]), .co(carry9[12]));
FA fa9_13(.a(sum8[14]), .b(A[13] & B[9]), .ci(carry9[12]), .s(sum9[13]), .co(carry9[13]));
FA fa9_14(.a(sum8[15]), .b(A[14] & B[9]), .ci(carry9[13]), .s(sum9[14]), .co(carry9[14]));
FA fa9_15(.a(sum8[16]), .b(A[15] & B[9]), .ci(carry9[14]), .s(sum9[15]), .co(carry9[15]));
FA fa9_16(.a(sum8[17]), .b(A[16] & B[9]), .ci(carry9[15]), .s(sum9[16]), .co(carry9[16]));
FA fa9_17(.a(sum8[18]), .b(A[17] & B[9]), .ci(carry9[16]), .s(sum9[17]), .co(carry9[17]));
FA fa9_18(.a(sum8[19]), .b(A[18] & B[9]), .ci(carry9[17]), .s(sum9[18]), .co(carry9[18]));
FA fa9_19(.a(sum8[20]), .b(A[19] & B[9]), .ci(carry9[18]), .s(sum9[19]), .co(carry9[19]));
FA fa9_20(.a(sum8[21]), .b(A[20] & B[9]), .ci(carry9[19]), .s(sum9[20]), .co(carry9[20]));
FA fa9_21(.a(sum8[22]), .b(A[21] & B[9]), .ci(carry9[20]), .s(sum9[21]), .co(carry9[21]));
FA fa9_22(.a(sum8[23]), .b(A[22] & B[9]), .ci(carry9[21]), .s(sum9[22]), .co(carry9[22]));
FA fa9_23(.a(sum8[24]), .b(A[23] & B[9]), .ci(carry9[22]), .s(sum9[23]), .co(carry9[23]));
FA fa9_24(.a(sum8[25]), .b(A[24] & B[9]), .ci(carry9[23]), .s(sum9[24]), .co(carry9[24]));
FA fa9_25(.a(sum8[26]), .b(A[25] & B[9]), .ci(carry9[24]), .s(sum9[25]), .co(carry9[25]));
FA fa9_26(.a(sum8[27]), .b(A[26] & B[9]), .ci(carry9[25]), .s(sum9[26]), .co(carry9[26]));
FA fa9_27(.a(sum8[28]), .b(A[27] & B[9]), .ci(carry9[26]), .s(sum9[27]), .co(carry9[27]));
FA fa9_28(.a(sum8[29]), .b(A[28] & B[9]), .ci(carry9[27]), .s(sum9[28]), .co(carry9[28]));
FA fa9_29(.a(sum8[30]), .b(A[29] & B[9]), .ci(carry9[28]), .s(sum9[29]), .co(carry9[29]));
FA fa9_30(.a(sum8[31]), .b(A[30] & B[9]), .ci(carry9[29]), .s(sum9[30]), .co(carry9[30]));
FA fa9_31(.a(carry8[31]), .b(A[31] & B[9]), .ci(carry9[30]), .s(sum9[31]), .co(carry9[31]));
FA fa10_0(.a(sum9[1]), .b(A[0] & B[10]), .ci(1'b0), .s(Z[10]), .co(carry10[0]));
FA fa10_1(.a(sum9[2]), .b(A[1] & B[10]), .ci(carry10[0]), .s(sum10[1]), .co(carry10[1]));
FA fa10_2(.a(sum9[3]), .b(A[2] & B[10]), .ci(carry10[1]), .s(sum10[2]), .co(carry10[2]));
FA fa10_3(.a(sum9[4]), .b(A[3] & B[10]), .ci(carry10[2]), .s(sum10[3]), .co(carry10[3]));
FA fa10_4(.a(sum9[5]), .b(A[4] & B[10]), .ci(carry10[3]), .s(sum10[4]), .co(carry10[4]));
FA fa10_5(.a(sum9[6]), .b(A[5] & B[10]), .ci(carry10[4]), .s(sum10[5]), .co(carry10[5]));
FA fa10_6(.a(sum9[7]), .b(A[6] & B[10]), .ci(carry10[5]), .s(sum10[6]), .co(carry10[6]));
FA fa10_7(.a(sum9[8]), .b(A[7] & B[10]), .ci(carry10[6]), .s(sum10[7]), .co(carry10[7]));
FA fa10_8(.a(sum9[9]), .b(A[8] & B[10]), .ci(carry10[7]), .s(sum10[8]), .co(carry10[8]));
FA fa10_9(.a(sum9[10]), .b(A[9] & B[10]), .ci(carry10[8]), .s(sum10[9]), .co(carry10[9]));
FA fa10_10(.a(sum9[11]), .b(A[10] & B[10]), .ci(carry10[9]), .s(sum10[10]), .co(carry10[10]));
FA fa10_11(.a(sum9[12]), .b(A[11] & B[10]), .ci(carry10[10]), .s(sum10[11]), .co(carry10[11]));
FA fa10_12(.a(sum9[13]), .b(A[12] & B[10]), .ci(carry10[11]), .s(sum10[12]), .co(carry10[12]));
FA fa10_13(.a(sum9[14]), .b(A[13] & B[10]), .ci(carry10[12]), .s(sum10[13]), .co(carry10[13]));
FA fa10_14(.a(sum9[15]), .b(A[14] & B[10]), .ci(carry10[13]), .s(sum10[14]), .co(carry10[14]));
FA fa10_15(.a(sum9[16]), .b(A[15] & B[10]), .ci(carry10[14]), .s(sum10[15]), .co(carry10[15]));
FA fa10_16(.a(sum9[17]), .b(A[16] & B[10]), .ci(carry10[15]), .s(sum10[16]), .co(carry10[16]));
FA fa10_17(.a(sum9[18]), .b(A[17] & B[10]), .ci(carry10[16]), .s(sum10[17]), .co(carry10[17]));
FA fa10_18(.a(sum9[19]), .b(A[18] & B[10]), .ci(carry10[17]), .s(sum10[18]), .co(carry10[18]));
FA fa10_19(.a(sum9[20]), .b(A[19] & B[10]), .ci(carry10[18]), .s(sum10[19]), .co(carry10[19]));
FA fa10_20(.a(sum9[21]), .b(A[20] & B[10]), .ci(carry10[19]), .s(sum10[20]), .co(carry10[20]));
FA fa10_21(.a(sum9[22]), .b(A[21] & B[10]), .ci(carry10[20]), .s(sum10[21]), .co(carry10[21]));
FA fa10_22(.a(sum9[23]), .b(A[22] & B[10]), .ci(carry10[21]), .s(sum10[22]), .co(carry10[22]));
FA fa10_23(.a(sum9[24]), .b(A[23] & B[10]), .ci(carry10[22]), .s(sum10[23]), .co(carry10[23]));
FA fa10_24(.a(sum9[25]), .b(A[24] & B[10]), .ci(carry10[23]), .s(sum10[24]), .co(carry10[24]));
FA fa10_25(.a(sum9[26]), .b(A[25] & B[10]), .ci(carry10[24]), .s(sum10[25]), .co(carry10[25]));
FA fa10_26(.a(sum9[27]), .b(A[26] & B[10]), .ci(carry10[25]), .s(sum10[26]), .co(carry10[26]));
FA fa10_27(.a(sum9[28]), .b(A[27] & B[10]), .ci(carry10[26]), .s(sum10[27]), .co(carry10[27]));
FA fa10_28(.a(sum9[29]), .b(A[28] & B[10]), .ci(carry10[27]), .s(sum10[28]), .co(carry10[28]));
FA fa10_29(.a(sum9[30]), .b(A[29] & B[10]), .ci(carry10[28]), .s(sum10[29]), .co(carry10[29]));
FA fa10_30(.a(sum9[31]), .b(A[30] & B[10]), .ci(carry10[29]), .s(sum10[30]), .co(carry10[30]));
FA fa10_31(.a(carry9[31]), .b(A[31] & B[10]), .ci(carry10[30]), .s(sum10[31]), .co(carry10[31]));
FA fa11_0(.a(sum10[1]), .b(A[0] & B[11]), .ci(1'b0), .s(Z[11]), .co(carry11[0]));
FA fa11_1(.a(sum10[2]), .b(A[1] & B[11]), .ci(carry11[0]), .s(sum11[1]), .co(carry11[1]));
FA fa11_2(.a(sum10[3]), .b(A[2] & B[11]), .ci(carry11[1]), .s(sum11[2]), .co(carry11[2]));
FA fa11_3(.a(sum10[4]), .b(A[3] & B[11]), .ci(carry11[2]), .s(sum11[3]), .co(carry11[3]));
FA fa11_4(.a(sum10[5]), .b(A[4] & B[11]), .ci(carry11[3]), .s(sum11[4]), .co(carry11[4]));
FA fa11_5(.a(sum10[6]), .b(A[5] & B[11]), .ci(carry11[4]), .s(sum11[5]), .co(carry11[5]));
FA fa11_6(.a(sum10[7]), .b(A[6] & B[11]), .ci(carry11[5]), .s(sum11[6]), .co(carry11[6]));
FA fa11_7(.a(sum10[8]), .b(A[7] & B[11]), .ci(carry11[6]), .s(sum11[7]), .co(carry11[7]));
FA fa11_8(.a(sum10[9]), .b(A[8] & B[11]), .ci(carry11[7]), .s(sum11[8]), .co(carry11[8]));
FA fa11_9(.a(sum10[10]), .b(A[9] & B[11]), .ci(carry11[8]), .s(sum11[9]), .co(carry11[9]));
FA fa11_10(.a(sum10[11]), .b(A[10] & B[11]), .ci(carry11[9]), .s(sum11[10]), .co(carry11[10]));
FA fa11_11(.a(sum10[12]), .b(A[11] & B[11]), .ci(carry11[10]), .s(sum11[11]), .co(carry11[11]));
FA fa11_12(.a(sum10[13]), .b(A[12] & B[11]), .ci(carry11[11]), .s(sum11[12]), .co(carry11[12]));
FA fa11_13(.a(sum10[14]), .b(A[13] & B[11]), .ci(carry11[12]), .s(sum11[13]), .co(carry11[13]));
FA fa11_14(.a(sum10[15]), .b(A[14] & B[11]), .ci(carry11[13]), .s(sum11[14]), .co(carry11[14]));
FA fa11_15(.a(sum10[16]), .b(A[15] & B[11]), .ci(carry11[14]), .s(sum11[15]), .co(carry11[15]));
FA fa11_16(.a(sum10[17]), .b(A[16] & B[11]), .ci(carry11[15]), .s(sum11[16]), .co(carry11[16]));
FA fa11_17(.a(sum10[18]), .b(A[17] & B[11]), .ci(carry11[16]), .s(sum11[17]), .co(carry11[17]));
FA fa11_18(.a(sum10[19]), .b(A[18] & B[11]), .ci(carry11[17]), .s(sum11[18]), .co(carry11[18]));
FA fa11_19(.a(sum10[20]), .b(A[19] & B[11]), .ci(carry11[18]), .s(sum11[19]), .co(carry11[19]));
FA fa11_20(.a(sum10[21]), .b(A[20] & B[11]), .ci(carry11[19]), .s(sum11[20]), .co(carry11[20]));
FA fa11_21(.a(sum10[22]), .b(A[21] & B[11]), .ci(carry11[20]), .s(sum11[21]), .co(carry11[21]));
FA fa11_22(.a(sum10[23]), .b(A[22] & B[11]), .ci(carry11[21]), .s(sum11[22]), .co(carry11[22]));
FA fa11_23(.a(sum10[24]), .b(A[23] & B[11]), .ci(carry11[22]), .s(sum11[23]), .co(carry11[23]));
FA fa11_24(.a(sum10[25]), .b(A[24] & B[11]), .ci(carry11[23]), .s(sum11[24]), .co(carry11[24]));
FA fa11_25(.a(sum10[26]), .b(A[25] & B[11]), .ci(carry11[24]), .s(sum11[25]), .co(carry11[25]));
FA fa11_26(.a(sum10[27]), .b(A[26] & B[11]), .ci(carry11[25]), .s(sum11[26]), .co(carry11[26]));
FA fa11_27(.a(sum10[28]), .b(A[27] & B[11]), .ci(carry11[26]), .s(sum11[27]), .co(carry11[27]));
FA fa11_28(.a(sum10[29]), .b(A[28] & B[11]), .ci(carry11[27]), .s(sum11[28]), .co(carry11[28]));
FA fa11_29(.a(sum10[30]), .b(A[29] & B[11]), .ci(carry11[28]), .s(sum11[29]), .co(carry11[29]));
FA fa11_30(.a(sum10[31]), .b(A[30] & B[11]), .ci(carry11[29]), .s(sum11[30]), .co(carry11[30]));
FA fa11_31(.a(carry10[31]), .b(A[31] & B[11]), .ci(carry11[30]), .s(sum11[31]), .co(carry11[31]));
FA fa12_0(.a(sum11[1]), .b(A[0] & B[12]), .ci(1'b0), .s(Z[12]), .co(carry12[0]));
FA fa12_1(.a(sum11[2]), .b(A[1] & B[12]), .ci(carry12[0]), .s(sum12[1]), .co(carry12[1]));
FA fa12_2(.a(sum11[3]), .b(A[2] & B[12]), .ci(carry12[1]), .s(sum12[2]), .co(carry12[2]));
FA fa12_3(.a(sum11[4]), .b(A[3] & B[12]), .ci(carry12[2]), .s(sum12[3]), .co(carry12[3]));
FA fa12_4(.a(sum11[5]), .b(A[4] & B[12]), .ci(carry12[3]), .s(sum12[4]), .co(carry12[4]));
FA fa12_5(.a(sum11[6]), .b(A[5] & B[12]), .ci(carry12[4]), .s(sum12[5]), .co(carry12[5]));
FA fa12_6(.a(sum11[7]), .b(A[6] & B[12]), .ci(carry12[5]), .s(sum12[6]), .co(carry12[6]));
FA fa12_7(.a(sum11[8]), .b(A[7] & B[12]), .ci(carry12[6]), .s(sum12[7]), .co(carry12[7]));
FA fa12_8(.a(sum11[9]), .b(A[8] & B[12]), .ci(carry12[7]), .s(sum12[8]), .co(carry12[8]));
FA fa12_9(.a(sum11[10]), .b(A[9] & B[12]), .ci(carry12[8]), .s(sum12[9]), .co(carry12[9]));
FA fa12_10(.a(sum11[11]), .b(A[10] & B[12]), .ci(carry12[9]), .s(sum12[10]), .co(carry12[10]));
FA fa12_11(.a(sum11[12]), .b(A[11] & B[12]), .ci(carry12[10]), .s(sum12[11]), .co(carry12[11]));
FA fa12_12(.a(sum11[13]), .b(A[12] & B[12]), .ci(carry12[11]), .s(sum12[12]), .co(carry12[12]));
FA fa12_13(.a(sum11[14]), .b(A[13] & B[12]), .ci(carry12[12]), .s(sum12[13]), .co(carry12[13]));
FA fa12_14(.a(sum11[15]), .b(A[14] & B[12]), .ci(carry12[13]), .s(sum12[14]), .co(carry12[14]));
FA fa12_15(.a(sum11[16]), .b(A[15] & B[12]), .ci(carry12[14]), .s(sum12[15]), .co(carry12[15]));
FA fa12_16(.a(sum11[17]), .b(A[16] & B[12]), .ci(carry12[15]), .s(sum12[16]), .co(carry12[16]));
FA fa12_17(.a(sum11[18]), .b(A[17] & B[12]), .ci(carry12[16]), .s(sum12[17]), .co(carry12[17]));
FA fa12_18(.a(sum11[19]), .b(A[18] & B[12]), .ci(carry12[17]), .s(sum12[18]), .co(carry12[18]));
FA fa12_19(.a(sum11[20]), .b(A[19] & B[12]), .ci(carry12[18]), .s(sum12[19]), .co(carry12[19]));
FA fa12_20(.a(sum11[21]), .b(A[20] & B[12]), .ci(carry12[19]), .s(sum12[20]), .co(carry12[20]));
FA fa12_21(.a(sum11[22]), .b(A[21] & B[12]), .ci(carry12[20]), .s(sum12[21]), .co(carry12[21]));
FA fa12_22(.a(sum11[23]), .b(A[22] & B[12]), .ci(carry12[21]), .s(sum12[22]), .co(carry12[22]));
FA fa12_23(.a(sum11[24]), .b(A[23] & B[12]), .ci(carry12[22]), .s(sum12[23]), .co(carry12[23]));
FA fa12_24(.a(sum11[25]), .b(A[24] & B[12]), .ci(carry12[23]), .s(sum12[24]), .co(carry12[24]));
FA fa12_25(.a(sum11[26]), .b(A[25] & B[12]), .ci(carry12[24]), .s(sum12[25]), .co(carry12[25]));
FA fa12_26(.a(sum11[27]), .b(A[26] & B[12]), .ci(carry12[25]), .s(sum12[26]), .co(carry12[26]));
FA fa12_27(.a(sum11[28]), .b(A[27] & B[12]), .ci(carry12[26]), .s(sum12[27]), .co(carry12[27]));
FA fa12_28(.a(sum11[29]), .b(A[28] & B[12]), .ci(carry12[27]), .s(sum12[28]), .co(carry12[28]));
FA fa12_29(.a(sum11[30]), .b(A[29] & B[12]), .ci(carry12[28]), .s(sum12[29]), .co(carry12[29]));
FA fa12_30(.a(sum11[31]), .b(A[30] & B[12]), .ci(carry12[29]), .s(sum12[30]), .co(carry12[30]));
FA fa12_31(.a(carry11[31]), .b(A[31] & B[12]), .ci(carry12[30]), .s(sum12[31]), .co(carry12[31]));
FA fa13_0(.a(sum12[1]), .b(A[0] & B[13]), .ci(1'b0), .s(Z[13]), .co(carry13[0]));
FA fa13_1(.a(sum12[2]), .b(A[1] & B[13]), .ci(carry13[0]), .s(sum13[1]), .co(carry13[1]));
FA fa13_2(.a(sum12[3]), .b(A[2] & B[13]), .ci(carry13[1]), .s(sum13[2]), .co(carry13[2]));
FA fa13_3(.a(sum12[4]), .b(A[3] & B[13]), .ci(carry13[2]), .s(sum13[3]), .co(carry13[3]));
FA fa13_4(.a(sum12[5]), .b(A[4] & B[13]), .ci(carry13[3]), .s(sum13[4]), .co(carry13[4]));
FA fa13_5(.a(sum12[6]), .b(A[5] & B[13]), .ci(carry13[4]), .s(sum13[5]), .co(carry13[5]));
FA fa13_6(.a(sum12[7]), .b(A[6] & B[13]), .ci(carry13[5]), .s(sum13[6]), .co(carry13[6]));
FA fa13_7(.a(sum12[8]), .b(A[7] & B[13]), .ci(carry13[6]), .s(sum13[7]), .co(carry13[7]));
FA fa13_8(.a(sum12[9]), .b(A[8] & B[13]), .ci(carry13[7]), .s(sum13[8]), .co(carry13[8]));
FA fa13_9(.a(sum12[10]), .b(A[9] & B[13]), .ci(carry13[8]), .s(sum13[9]), .co(carry13[9]));
FA fa13_10(.a(sum12[11]), .b(A[10] & B[13]), .ci(carry13[9]), .s(sum13[10]), .co(carry13[10]));
FA fa13_11(.a(sum12[12]), .b(A[11] & B[13]), .ci(carry13[10]), .s(sum13[11]), .co(carry13[11]));
FA fa13_12(.a(sum12[13]), .b(A[12] & B[13]), .ci(carry13[11]), .s(sum13[12]), .co(carry13[12]));
FA fa13_13(.a(sum12[14]), .b(A[13] & B[13]), .ci(carry13[12]), .s(sum13[13]), .co(carry13[13]));
FA fa13_14(.a(sum12[15]), .b(A[14] & B[13]), .ci(carry13[13]), .s(sum13[14]), .co(carry13[14]));
FA fa13_15(.a(sum12[16]), .b(A[15] & B[13]), .ci(carry13[14]), .s(sum13[15]), .co(carry13[15]));
FA fa13_16(.a(sum12[17]), .b(A[16] & B[13]), .ci(carry13[15]), .s(sum13[16]), .co(carry13[16]));
FA fa13_17(.a(sum12[18]), .b(A[17] & B[13]), .ci(carry13[16]), .s(sum13[17]), .co(carry13[17]));
FA fa13_18(.a(sum12[19]), .b(A[18] & B[13]), .ci(carry13[17]), .s(sum13[18]), .co(carry13[18]));
FA fa13_19(.a(sum12[20]), .b(A[19] & B[13]), .ci(carry13[18]), .s(sum13[19]), .co(carry13[19]));
FA fa13_20(.a(sum12[21]), .b(A[20] & B[13]), .ci(carry13[19]), .s(sum13[20]), .co(carry13[20]));
FA fa13_21(.a(sum12[22]), .b(A[21] & B[13]), .ci(carry13[20]), .s(sum13[21]), .co(carry13[21]));
FA fa13_22(.a(sum12[23]), .b(A[22] & B[13]), .ci(carry13[21]), .s(sum13[22]), .co(carry13[22]));
FA fa13_23(.a(sum12[24]), .b(A[23] & B[13]), .ci(carry13[22]), .s(sum13[23]), .co(carry13[23]));
FA fa13_24(.a(sum12[25]), .b(A[24] & B[13]), .ci(carry13[23]), .s(sum13[24]), .co(carry13[24]));
FA fa13_25(.a(sum12[26]), .b(A[25] & B[13]), .ci(carry13[24]), .s(sum13[25]), .co(carry13[25]));
FA fa13_26(.a(sum12[27]), .b(A[26] & B[13]), .ci(carry13[25]), .s(sum13[26]), .co(carry13[26]));
FA fa13_27(.a(sum12[28]), .b(A[27] & B[13]), .ci(carry13[26]), .s(sum13[27]), .co(carry13[27]));
FA fa13_28(.a(sum12[29]), .b(A[28] & B[13]), .ci(carry13[27]), .s(sum13[28]), .co(carry13[28]));
FA fa13_29(.a(sum12[30]), .b(A[29] & B[13]), .ci(carry13[28]), .s(sum13[29]), .co(carry13[29]));
FA fa13_30(.a(sum12[31]), .b(A[30] & B[13]), .ci(carry13[29]), .s(sum13[30]), .co(carry13[30]));
FA fa13_31(.a(carry12[31]), .b(A[31] & B[13]), .ci(carry13[30]), .s(sum13[31]), .co(carry13[31]));
FA fa14_0(.a(sum13[1]), .b(A[0] & B[14]), .ci(1'b0), .s(Z[14]), .co(carry14[0]));
FA fa14_1(.a(sum13[2]), .b(A[1] & B[14]), .ci(carry14[0]), .s(sum14[1]), .co(carry14[1]));
FA fa14_2(.a(sum13[3]), .b(A[2] & B[14]), .ci(carry14[1]), .s(sum14[2]), .co(carry14[2]));
FA fa14_3(.a(sum13[4]), .b(A[3] & B[14]), .ci(carry14[2]), .s(sum14[3]), .co(carry14[3]));
FA fa14_4(.a(sum13[5]), .b(A[4] & B[14]), .ci(carry14[3]), .s(sum14[4]), .co(carry14[4]));
FA fa14_5(.a(sum13[6]), .b(A[5] & B[14]), .ci(carry14[4]), .s(sum14[5]), .co(carry14[5]));
FA fa14_6(.a(sum13[7]), .b(A[6] & B[14]), .ci(carry14[5]), .s(sum14[6]), .co(carry14[6]));
FA fa14_7(.a(sum13[8]), .b(A[7] & B[14]), .ci(carry14[6]), .s(sum14[7]), .co(carry14[7]));
FA fa14_8(.a(sum13[9]), .b(A[8] & B[14]), .ci(carry14[7]), .s(sum14[8]), .co(carry14[8]));
FA fa14_9(.a(sum13[10]), .b(A[9] & B[14]), .ci(carry14[8]), .s(sum14[9]), .co(carry14[9]));
FA fa14_10(.a(sum13[11]), .b(A[10] & B[14]), .ci(carry14[9]), .s(sum14[10]), .co(carry14[10]));
FA fa14_11(.a(sum13[12]), .b(A[11] & B[14]), .ci(carry14[10]), .s(sum14[11]), .co(carry14[11]));
FA fa14_12(.a(sum13[13]), .b(A[12] & B[14]), .ci(carry14[11]), .s(sum14[12]), .co(carry14[12]));
FA fa14_13(.a(sum13[14]), .b(A[13] & B[14]), .ci(carry14[12]), .s(sum14[13]), .co(carry14[13]));
FA fa14_14(.a(sum13[15]), .b(A[14] & B[14]), .ci(carry14[13]), .s(sum14[14]), .co(carry14[14]));
FA fa14_15(.a(sum13[16]), .b(A[15] & B[14]), .ci(carry14[14]), .s(sum14[15]), .co(carry14[15]));
FA fa14_16(.a(sum13[17]), .b(A[16] & B[14]), .ci(carry14[15]), .s(sum14[16]), .co(carry14[16]));
FA fa14_17(.a(sum13[18]), .b(A[17] & B[14]), .ci(carry14[16]), .s(sum14[17]), .co(carry14[17]));
FA fa14_18(.a(sum13[19]), .b(A[18] & B[14]), .ci(carry14[17]), .s(sum14[18]), .co(carry14[18]));
FA fa14_19(.a(sum13[20]), .b(A[19] & B[14]), .ci(carry14[18]), .s(sum14[19]), .co(carry14[19]));
FA fa14_20(.a(sum13[21]), .b(A[20] & B[14]), .ci(carry14[19]), .s(sum14[20]), .co(carry14[20]));
FA fa14_21(.a(sum13[22]), .b(A[21] & B[14]), .ci(carry14[20]), .s(sum14[21]), .co(carry14[21]));
FA fa14_22(.a(sum13[23]), .b(A[22] & B[14]), .ci(carry14[21]), .s(sum14[22]), .co(carry14[22]));
FA fa14_23(.a(sum13[24]), .b(A[23] & B[14]), .ci(carry14[22]), .s(sum14[23]), .co(carry14[23]));
FA fa14_24(.a(sum13[25]), .b(A[24] & B[14]), .ci(carry14[23]), .s(sum14[24]), .co(carry14[24]));
FA fa14_25(.a(sum13[26]), .b(A[25] & B[14]), .ci(carry14[24]), .s(sum14[25]), .co(carry14[25]));
FA fa14_26(.a(sum13[27]), .b(A[26] & B[14]), .ci(carry14[25]), .s(sum14[26]), .co(carry14[26]));
FA fa14_27(.a(sum13[28]), .b(A[27] & B[14]), .ci(carry14[26]), .s(sum14[27]), .co(carry14[27]));
FA fa14_28(.a(sum13[29]), .b(A[28] & B[14]), .ci(carry14[27]), .s(sum14[28]), .co(carry14[28]));
FA fa14_29(.a(sum13[30]), .b(A[29] & B[14]), .ci(carry14[28]), .s(sum14[29]), .co(carry14[29]));
FA fa14_30(.a(sum13[31]), .b(A[30] & B[14]), .ci(carry14[29]), .s(sum14[30]), .co(carry14[30]));
FA fa14_31(.a(carry13[31]), .b(A[31] & B[14]), .ci(carry14[30]), .s(sum14[31]), .co(carry14[31]));
FA fa15_0(.a(sum14[1]), .b(A[0] & B[15]), .ci(1'b0), .s(Z[15]), .co(carry15[0]));
FA fa15_1(.a(sum14[2]), .b(A[1] & B[15]), .ci(carry15[0]), .s(sum15[1]), .co(carry15[1]));
FA fa15_2(.a(sum14[3]), .b(A[2] & B[15]), .ci(carry15[1]), .s(sum15[2]), .co(carry15[2]));
FA fa15_3(.a(sum14[4]), .b(A[3] & B[15]), .ci(carry15[2]), .s(sum15[3]), .co(carry15[3]));
FA fa15_4(.a(sum14[5]), .b(A[4] & B[15]), .ci(carry15[3]), .s(sum15[4]), .co(carry15[4]));
FA fa15_5(.a(sum14[6]), .b(A[5] & B[15]), .ci(carry15[4]), .s(sum15[5]), .co(carry15[5]));
FA fa15_6(.a(sum14[7]), .b(A[6] & B[15]), .ci(carry15[5]), .s(sum15[6]), .co(carry15[6]));
FA fa15_7(.a(sum14[8]), .b(A[7] & B[15]), .ci(carry15[6]), .s(sum15[7]), .co(carry15[7]));
FA fa15_8(.a(sum14[9]), .b(A[8] & B[15]), .ci(carry15[7]), .s(sum15[8]), .co(carry15[8]));
FA fa15_9(.a(sum14[10]), .b(A[9] & B[15]), .ci(carry15[8]), .s(sum15[9]), .co(carry15[9]));
FA fa15_10(.a(sum14[11]), .b(A[10] & B[15]), .ci(carry15[9]), .s(sum15[10]), .co(carry15[10]));
FA fa15_11(.a(sum14[12]), .b(A[11] & B[15]), .ci(carry15[10]), .s(sum15[11]), .co(carry15[11]));
FA fa15_12(.a(sum14[13]), .b(A[12] & B[15]), .ci(carry15[11]), .s(sum15[12]), .co(carry15[12]));
FA fa15_13(.a(sum14[14]), .b(A[13] & B[15]), .ci(carry15[12]), .s(sum15[13]), .co(carry15[13]));
FA fa15_14(.a(sum14[15]), .b(A[14] & B[15]), .ci(carry15[13]), .s(sum15[14]), .co(carry15[14]));
FA fa15_15(.a(sum14[16]), .b(A[15] & B[15]), .ci(carry15[14]), .s(sum15[15]), .co(carry15[15]));
FA fa15_16(.a(sum14[17]), .b(A[16] & B[15]), .ci(carry15[15]), .s(sum15[16]), .co(carry15[16]));
FA fa15_17(.a(sum14[18]), .b(A[17] & B[15]), .ci(carry15[16]), .s(sum15[17]), .co(carry15[17]));
FA fa15_18(.a(sum14[19]), .b(A[18] & B[15]), .ci(carry15[17]), .s(sum15[18]), .co(carry15[18]));
FA fa15_19(.a(sum14[20]), .b(A[19] & B[15]), .ci(carry15[18]), .s(sum15[19]), .co(carry15[19]));
FA fa15_20(.a(sum14[21]), .b(A[20] & B[15]), .ci(carry15[19]), .s(sum15[20]), .co(carry15[20]));
FA fa15_21(.a(sum14[22]), .b(A[21] & B[15]), .ci(carry15[20]), .s(sum15[21]), .co(carry15[21]));
FA fa15_22(.a(sum14[23]), .b(A[22] & B[15]), .ci(carry15[21]), .s(sum15[22]), .co(carry15[22]));
FA fa15_23(.a(sum14[24]), .b(A[23] & B[15]), .ci(carry15[22]), .s(sum15[23]), .co(carry15[23]));
FA fa15_24(.a(sum14[25]), .b(A[24] & B[15]), .ci(carry15[23]), .s(sum15[24]), .co(carry15[24]));
FA fa15_25(.a(sum14[26]), .b(A[25] & B[15]), .ci(carry15[24]), .s(sum15[25]), .co(carry15[25]));
FA fa15_26(.a(sum14[27]), .b(A[26] & B[15]), .ci(carry15[25]), .s(sum15[26]), .co(carry15[26]));
FA fa15_27(.a(sum14[28]), .b(A[27] & B[15]), .ci(carry15[26]), .s(sum15[27]), .co(carry15[27]));
FA fa15_28(.a(sum14[29]), .b(A[28] & B[15]), .ci(carry15[27]), .s(sum15[28]), .co(carry15[28]));
FA fa15_29(.a(sum14[30]), .b(A[29] & B[15]), .ci(carry15[28]), .s(sum15[29]), .co(carry15[29]));
FA fa15_30(.a(sum14[31]), .b(A[30] & B[15]), .ci(carry15[29]), .s(sum15[30]), .co(carry15[30]));
FA fa15_31(.a(carry14[31]), .b(A[31] & B[15]), .ci(carry15[30]), .s(sum15[31]), .co(carry15[31]));
FA fa16_0(.a(sum15[1]), .b(A[0] & B[16]), .ci(1'b0), .s(Z[16]), .co(carry16[0]));
FA fa16_1(.a(sum15[2]), .b(A[1] & B[16]), .ci(carry16[0]), .s(sum16[1]), .co(carry16[1]));
FA fa16_2(.a(sum15[3]), .b(A[2] & B[16]), .ci(carry16[1]), .s(sum16[2]), .co(carry16[2]));
FA fa16_3(.a(sum15[4]), .b(A[3] & B[16]), .ci(carry16[2]), .s(sum16[3]), .co(carry16[3]));
FA fa16_4(.a(sum15[5]), .b(A[4] & B[16]), .ci(carry16[3]), .s(sum16[4]), .co(carry16[4]));
FA fa16_5(.a(sum15[6]), .b(A[5] & B[16]), .ci(carry16[4]), .s(sum16[5]), .co(carry16[5]));
FA fa16_6(.a(sum15[7]), .b(A[6] & B[16]), .ci(carry16[5]), .s(sum16[6]), .co(carry16[6]));
FA fa16_7(.a(sum15[8]), .b(A[7] & B[16]), .ci(carry16[6]), .s(sum16[7]), .co(carry16[7]));
FA fa16_8(.a(sum15[9]), .b(A[8] & B[16]), .ci(carry16[7]), .s(sum16[8]), .co(carry16[8]));
FA fa16_9(.a(sum15[10]), .b(A[9] & B[16]), .ci(carry16[8]), .s(sum16[9]), .co(carry16[9]));
FA fa16_10(.a(sum15[11]), .b(A[10] & B[16]), .ci(carry16[9]), .s(sum16[10]), .co(carry16[10]));
FA fa16_11(.a(sum15[12]), .b(A[11] & B[16]), .ci(carry16[10]), .s(sum16[11]), .co(carry16[11]));
FA fa16_12(.a(sum15[13]), .b(A[12] & B[16]), .ci(carry16[11]), .s(sum16[12]), .co(carry16[12]));
FA fa16_13(.a(sum15[14]), .b(A[13] & B[16]), .ci(carry16[12]), .s(sum16[13]), .co(carry16[13]));
FA fa16_14(.a(sum15[15]), .b(A[14] & B[16]), .ci(carry16[13]), .s(sum16[14]), .co(carry16[14]));
FA fa16_15(.a(sum15[16]), .b(A[15] & B[16]), .ci(carry16[14]), .s(sum16[15]), .co(carry16[15]));
FA fa16_16(.a(sum15[17]), .b(A[16] & B[16]), .ci(carry16[15]), .s(sum16[16]), .co(carry16[16]));
FA fa16_17(.a(sum15[18]), .b(A[17] & B[16]), .ci(carry16[16]), .s(sum16[17]), .co(carry16[17]));
FA fa16_18(.a(sum15[19]), .b(A[18] & B[16]), .ci(carry16[17]), .s(sum16[18]), .co(carry16[18]));
FA fa16_19(.a(sum15[20]), .b(A[19] & B[16]), .ci(carry16[18]), .s(sum16[19]), .co(carry16[19]));
FA fa16_20(.a(sum15[21]), .b(A[20] & B[16]), .ci(carry16[19]), .s(sum16[20]), .co(carry16[20]));
FA fa16_21(.a(sum15[22]), .b(A[21] & B[16]), .ci(carry16[20]), .s(sum16[21]), .co(carry16[21]));
FA fa16_22(.a(sum15[23]), .b(A[22] & B[16]), .ci(carry16[21]), .s(sum16[22]), .co(carry16[22]));
FA fa16_23(.a(sum15[24]), .b(A[23] & B[16]), .ci(carry16[22]), .s(sum16[23]), .co(carry16[23]));
FA fa16_24(.a(sum15[25]), .b(A[24] & B[16]), .ci(carry16[23]), .s(sum16[24]), .co(carry16[24]));
FA fa16_25(.a(sum15[26]), .b(A[25] & B[16]), .ci(carry16[24]), .s(sum16[25]), .co(carry16[25]));
FA fa16_26(.a(sum15[27]), .b(A[26] & B[16]), .ci(carry16[25]), .s(sum16[26]), .co(carry16[26]));
FA fa16_27(.a(sum15[28]), .b(A[27] & B[16]), .ci(carry16[26]), .s(sum16[27]), .co(carry16[27]));
FA fa16_28(.a(sum15[29]), .b(A[28] & B[16]), .ci(carry16[27]), .s(sum16[28]), .co(carry16[28]));
FA fa16_29(.a(sum15[30]), .b(A[29] & B[16]), .ci(carry16[28]), .s(sum16[29]), .co(carry16[29]));
FA fa16_30(.a(sum15[31]), .b(A[30] & B[16]), .ci(carry16[29]), .s(sum16[30]), .co(carry16[30]));
FA fa16_31(.a(carry15[31]), .b(A[31] & B[16]), .ci(carry16[30]), .s(sum16[31]), .co(carry16[31]));
FA fa17_0(.a(sum16[1]), .b(A[0] & B[17]), .ci(1'b0), .s(Z[17]), .co(carry17[0]));
FA fa17_1(.a(sum16[2]), .b(A[1] & B[17]), .ci(carry17[0]), .s(sum17[1]), .co(carry17[1]));
FA fa17_2(.a(sum16[3]), .b(A[2] & B[17]), .ci(carry17[1]), .s(sum17[2]), .co(carry17[2]));
FA fa17_3(.a(sum16[4]), .b(A[3] & B[17]), .ci(carry17[2]), .s(sum17[3]), .co(carry17[3]));
FA fa17_4(.a(sum16[5]), .b(A[4] & B[17]), .ci(carry17[3]), .s(sum17[4]), .co(carry17[4]));
FA fa17_5(.a(sum16[6]), .b(A[5] & B[17]), .ci(carry17[4]), .s(sum17[5]), .co(carry17[5]));
FA fa17_6(.a(sum16[7]), .b(A[6] & B[17]), .ci(carry17[5]), .s(sum17[6]), .co(carry17[6]));
FA fa17_7(.a(sum16[8]), .b(A[7] & B[17]), .ci(carry17[6]), .s(sum17[7]), .co(carry17[7]));
FA fa17_8(.a(sum16[9]), .b(A[8] & B[17]), .ci(carry17[7]), .s(sum17[8]), .co(carry17[8]));
FA fa17_9(.a(sum16[10]), .b(A[9] & B[17]), .ci(carry17[8]), .s(sum17[9]), .co(carry17[9]));
FA fa17_10(.a(sum16[11]), .b(A[10] & B[17]), .ci(carry17[9]), .s(sum17[10]), .co(carry17[10]));
FA fa17_11(.a(sum16[12]), .b(A[11] & B[17]), .ci(carry17[10]), .s(sum17[11]), .co(carry17[11]));
FA fa17_12(.a(sum16[13]), .b(A[12] & B[17]), .ci(carry17[11]), .s(sum17[12]), .co(carry17[12]));
FA fa17_13(.a(sum16[14]), .b(A[13] & B[17]), .ci(carry17[12]), .s(sum17[13]), .co(carry17[13]));
FA fa17_14(.a(sum16[15]), .b(A[14] & B[17]), .ci(carry17[13]), .s(sum17[14]), .co(carry17[14]));
FA fa17_15(.a(sum16[16]), .b(A[15] & B[17]), .ci(carry17[14]), .s(sum17[15]), .co(carry17[15]));
FA fa17_16(.a(sum16[17]), .b(A[16] & B[17]), .ci(carry17[15]), .s(sum17[16]), .co(carry17[16]));
FA fa17_17(.a(sum16[18]), .b(A[17] & B[17]), .ci(carry17[16]), .s(sum17[17]), .co(carry17[17]));
FA fa17_18(.a(sum16[19]), .b(A[18] & B[17]), .ci(carry17[17]), .s(sum17[18]), .co(carry17[18]));
FA fa17_19(.a(sum16[20]), .b(A[19] & B[17]), .ci(carry17[18]), .s(sum17[19]), .co(carry17[19]));
FA fa17_20(.a(sum16[21]), .b(A[20] & B[17]), .ci(carry17[19]), .s(sum17[20]), .co(carry17[20]));
FA fa17_21(.a(sum16[22]), .b(A[21] & B[17]), .ci(carry17[20]), .s(sum17[21]), .co(carry17[21]));
FA fa17_22(.a(sum16[23]), .b(A[22] & B[17]), .ci(carry17[21]), .s(sum17[22]), .co(carry17[22]));
FA fa17_23(.a(sum16[24]), .b(A[23] & B[17]), .ci(carry17[22]), .s(sum17[23]), .co(carry17[23]));
FA fa17_24(.a(sum16[25]), .b(A[24] & B[17]), .ci(carry17[23]), .s(sum17[24]), .co(carry17[24]));
FA fa17_25(.a(sum16[26]), .b(A[25] & B[17]), .ci(carry17[24]), .s(sum17[25]), .co(carry17[25]));
FA fa17_26(.a(sum16[27]), .b(A[26] & B[17]), .ci(carry17[25]), .s(sum17[26]), .co(carry17[26]));
FA fa17_27(.a(sum16[28]), .b(A[27] & B[17]), .ci(carry17[26]), .s(sum17[27]), .co(carry17[27]));
FA fa17_28(.a(sum16[29]), .b(A[28] & B[17]), .ci(carry17[27]), .s(sum17[28]), .co(carry17[28]));
FA fa17_29(.a(sum16[30]), .b(A[29] & B[17]), .ci(carry17[28]), .s(sum17[29]), .co(carry17[29]));
FA fa17_30(.a(sum16[31]), .b(A[30] & B[17]), .ci(carry17[29]), .s(sum17[30]), .co(carry17[30]));
FA fa17_31(.a(carry16[31]), .b(A[31] & B[17]), .ci(carry17[30]), .s(sum17[31]), .co(carry17[31]));
FA fa18_0(.a(sum17[1]), .b(A[0] & B[18]), .ci(1'b0), .s(Z[18]), .co(carry18[0]));
FA fa18_1(.a(sum17[2]), .b(A[1] & B[18]), .ci(carry18[0]), .s(sum18[1]), .co(carry18[1]));
FA fa18_2(.a(sum17[3]), .b(A[2] & B[18]), .ci(carry18[1]), .s(sum18[2]), .co(carry18[2]));
FA fa18_3(.a(sum17[4]), .b(A[3] & B[18]), .ci(carry18[2]), .s(sum18[3]), .co(carry18[3]));
FA fa18_4(.a(sum17[5]), .b(A[4] & B[18]), .ci(carry18[3]), .s(sum18[4]), .co(carry18[4]));
FA fa18_5(.a(sum17[6]), .b(A[5] & B[18]), .ci(carry18[4]), .s(sum18[5]), .co(carry18[5]));
FA fa18_6(.a(sum17[7]), .b(A[6] & B[18]), .ci(carry18[5]), .s(sum18[6]), .co(carry18[6]));
FA fa18_7(.a(sum17[8]), .b(A[7] & B[18]), .ci(carry18[6]), .s(sum18[7]), .co(carry18[7]));
FA fa18_8(.a(sum17[9]), .b(A[8] & B[18]), .ci(carry18[7]), .s(sum18[8]), .co(carry18[8]));
FA fa18_9(.a(sum17[10]), .b(A[9] & B[18]), .ci(carry18[8]), .s(sum18[9]), .co(carry18[9]));
FA fa18_10(.a(sum17[11]), .b(A[10] & B[18]), .ci(carry18[9]), .s(sum18[10]), .co(carry18[10]));
FA fa18_11(.a(sum17[12]), .b(A[11] & B[18]), .ci(carry18[10]), .s(sum18[11]), .co(carry18[11]));
FA fa18_12(.a(sum17[13]), .b(A[12] & B[18]), .ci(carry18[11]), .s(sum18[12]), .co(carry18[12]));
FA fa18_13(.a(sum17[14]), .b(A[13] & B[18]), .ci(carry18[12]), .s(sum18[13]), .co(carry18[13]));
FA fa18_14(.a(sum17[15]), .b(A[14] & B[18]), .ci(carry18[13]), .s(sum18[14]), .co(carry18[14]));
FA fa18_15(.a(sum17[16]), .b(A[15] & B[18]), .ci(carry18[14]), .s(sum18[15]), .co(carry18[15]));
FA fa18_16(.a(sum17[17]), .b(A[16] & B[18]), .ci(carry18[15]), .s(sum18[16]), .co(carry18[16]));
FA fa18_17(.a(sum17[18]), .b(A[17] & B[18]), .ci(carry18[16]), .s(sum18[17]), .co(carry18[17]));
FA fa18_18(.a(sum17[19]), .b(A[18] & B[18]), .ci(carry18[17]), .s(sum18[18]), .co(carry18[18]));
FA fa18_19(.a(sum17[20]), .b(A[19] & B[18]), .ci(carry18[18]), .s(sum18[19]), .co(carry18[19]));
FA fa18_20(.a(sum17[21]), .b(A[20] & B[18]), .ci(carry18[19]), .s(sum18[20]), .co(carry18[20]));
FA fa18_21(.a(sum17[22]), .b(A[21] & B[18]), .ci(carry18[20]), .s(sum18[21]), .co(carry18[21]));
FA fa18_22(.a(sum17[23]), .b(A[22] & B[18]), .ci(carry18[21]), .s(sum18[22]), .co(carry18[22]));
FA fa18_23(.a(sum17[24]), .b(A[23] & B[18]), .ci(carry18[22]), .s(sum18[23]), .co(carry18[23]));
FA fa18_24(.a(sum17[25]), .b(A[24] & B[18]), .ci(carry18[23]), .s(sum18[24]), .co(carry18[24]));
FA fa18_25(.a(sum17[26]), .b(A[25] & B[18]), .ci(carry18[24]), .s(sum18[25]), .co(carry18[25]));
FA fa18_26(.a(sum17[27]), .b(A[26] & B[18]), .ci(carry18[25]), .s(sum18[26]), .co(carry18[26]));
FA fa18_27(.a(sum17[28]), .b(A[27] & B[18]), .ci(carry18[26]), .s(sum18[27]), .co(carry18[27]));
FA fa18_28(.a(sum17[29]), .b(A[28] & B[18]), .ci(carry18[27]), .s(sum18[28]), .co(carry18[28]));
FA fa18_29(.a(sum17[30]), .b(A[29] & B[18]), .ci(carry18[28]), .s(sum18[29]), .co(carry18[29]));
FA fa18_30(.a(sum17[31]), .b(A[30] & B[18]), .ci(carry18[29]), .s(sum18[30]), .co(carry18[30]));
FA fa18_31(.a(carry17[31]), .b(A[31] & B[18]), .ci(carry18[30]), .s(sum18[31]), .co(carry18[31]));
FA fa19_0(.a(sum18[1]), .b(A[0] & B[19]), .ci(1'b0), .s(Z[19]), .co(carry19[0]));
FA fa19_1(.a(sum18[2]), .b(A[1] & B[19]), .ci(carry19[0]), .s(sum19[1]), .co(carry19[1]));
FA fa19_2(.a(sum18[3]), .b(A[2] & B[19]), .ci(carry19[1]), .s(sum19[2]), .co(carry19[2]));
FA fa19_3(.a(sum18[4]), .b(A[3] & B[19]), .ci(carry19[2]), .s(sum19[3]), .co(carry19[3]));
FA fa19_4(.a(sum18[5]), .b(A[4] & B[19]), .ci(carry19[3]), .s(sum19[4]), .co(carry19[4]));
FA fa19_5(.a(sum18[6]), .b(A[5] & B[19]), .ci(carry19[4]), .s(sum19[5]), .co(carry19[5]));
FA fa19_6(.a(sum18[7]), .b(A[6] & B[19]), .ci(carry19[5]), .s(sum19[6]), .co(carry19[6]));
FA fa19_7(.a(sum18[8]), .b(A[7] & B[19]), .ci(carry19[6]), .s(sum19[7]), .co(carry19[7]));
FA fa19_8(.a(sum18[9]), .b(A[8] & B[19]), .ci(carry19[7]), .s(sum19[8]), .co(carry19[8]));
FA fa19_9(.a(sum18[10]), .b(A[9] & B[19]), .ci(carry19[8]), .s(sum19[9]), .co(carry19[9]));
FA fa19_10(.a(sum18[11]), .b(A[10] & B[19]), .ci(carry19[9]), .s(sum19[10]), .co(carry19[10]));
FA fa19_11(.a(sum18[12]), .b(A[11] & B[19]), .ci(carry19[10]), .s(sum19[11]), .co(carry19[11]));
FA fa19_12(.a(sum18[13]), .b(A[12] & B[19]), .ci(carry19[11]), .s(sum19[12]), .co(carry19[12]));
FA fa19_13(.a(sum18[14]), .b(A[13] & B[19]), .ci(carry19[12]), .s(sum19[13]), .co(carry19[13]));
FA fa19_14(.a(sum18[15]), .b(A[14] & B[19]), .ci(carry19[13]), .s(sum19[14]), .co(carry19[14]));
FA fa19_15(.a(sum18[16]), .b(A[15] & B[19]), .ci(carry19[14]), .s(sum19[15]), .co(carry19[15]));
FA fa19_16(.a(sum18[17]), .b(A[16] & B[19]), .ci(carry19[15]), .s(sum19[16]), .co(carry19[16]));
FA fa19_17(.a(sum18[18]), .b(A[17] & B[19]), .ci(carry19[16]), .s(sum19[17]), .co(carry19[17]));
FA fa19_18(.a(sum18[19]), .b(A[18] & B[19]), .ci(carry19[17]), .s(sum19[18]), .co(carry19[18]));
FA fa19_19(.a(sum18[20]), .b(A[19] & B[19]), .ci(carry19[18]), .s(sum19[19]), .co(carry19[19]));
FA fa19_20(.a(sum18[21]), .b(A[20] & B[19]), .ci(carry19[19]), .s(sum19[20]), .co(carry19[20]));
FA fa19_21(.a(sum18[22]), .b(A[21] & B[19]), .ci(carry19[20]), .s(sum19[21]), .co(carry19[21]));
FA fa19_22(.a(sum18[23]), .b(A[22] & B[19]), .ci(carry19[21]), .s(sum19[22]), .co(carry19[22]));
FA fa19_23(.a(sum18[24]), .b(A[23] & B[19]), .ci(carry19[22]), .s(sum19[23]), .co(carry19[23]));
FA fa19_24(.a(sum18[25]), .b(A[24] & B[19]), .ci(carry19[23]), .s(sum19[24]), .co(carry19[24]));
FA fa19_25(.a(sum18[26]), .b(A[25] & B[19]), .ci(carry19[24]), .s(sum19[25]), .co(carry19[25]));
FA fa19_26(.a(sum18[27]), .b(A[26] & B[19]), .ci(carry19[25]), .s(sum19[26]), .co(carry19[26]));
FA fa19_27(.a(sum18[28]), .b(A[27] & B[19]), .ci(carry19[26]), .s(sum19[27]), .co(carry19[27]));
FA fa19_28(.a(sum18[29]), .b(A[28] & B[19]), .ci(carry19[27]), .s(sum19[28]), .co(carry19[28]));
FA fa19_29(.a(sum18[30]), .b(A[29] & B[19]), .ci(carry19[28]), .s(sum19[29]), .co(carry19[29]));
FA fa19_30(.a(sum18[31]), .b(A[30] & B[19]), .ci(carry19[29]), .s(sum19[30]), .co(carry19[30]));
FA fa19_31(.a(carry18[31]), .b(A[31] & B[19]), .ci(carry19[30]), .s(sum19[31]), .co(carry19[31]));
FA fa20_0(.a(sum19[1]), .b(A[0] & B[20]), .ci(1'b0), .s(Z[20]), .co(carry20[0]));
FA fa20_1(.a(sum19[2]), .b(A[1] & B[20]), .ci(carry20[0]), .s(sum20[1]), .co(carry20[1]));
FA fa20_2(.a(sum19[3]), .b(A[2] & B[20]), .ci(carry20[1]), .s(sum20[2]), .co(carry20[2]));
FA fa20_3(.a(sum19[4]), .b(A[3] & B[20]), .ci(carry20[2]), .s(sum20[3]), .co(carry20[3]));
FA fa20_4(.a(sum19[5]), .b(A[4] & B[20]), .ci(carry20[3]), .s(sum20[4]), .co(carry20[4]));
FA fa20_5(.a(sum19[6]), .b(A[5] & B[20]), .ci(carry20[4]), .s(sum20[5]), .co(carry20[5]));
FA fa20_6(.a(sum19[7]), .b(A[6] & B[20]), .ci(carry20[5]), .s(sum20[6]), .co(carry20[6]));
FA fa20_7(.a(sum19[8]), .b(A[7] & B[20]), .ci(carry20[6]), .s(sum20[7]), .co(carry20[7]));
FA fa20_8(.a(sum19[9]), .b(A[8] & B[20]), .ci(carry20[7]), .s(sum20[8]), .co(carry20[8]));
FA fa20_9(.a(sum19[10]), .b(A[9] & B[20]), .ci(carry20[8]), .s(sum20[9]), .co(carry20[9]));
FA fa20_10(.a(sum19[11]), .b(A[10] & B[20]), .ci(carry20[9]), .s(sum20[10]), .co(carry20[10]));
FA fa20_11(.a(sum19[12]), .b(A[11] & B[20]), .ci(carry20[10]), .s(sum20[11]), .co(carry20[11]));
FA fa20_12(.a(sum19[13]), .b(A[12] & B[20]), .ci(carry20[11]), .s(sum20[12]), .co(carry20[12]));
FA fa20_13(.a(sum19[14]), .b(A[13] & B[20]), .ci(carry20[12]), .s(sum20[13]), .co(carry20[13]));
FA fa20_14(.a(sum19[15]), .b(A[14] & B[20]), .ci(carry20[13]), .s(sum20[14]), .co(carry20[14]));
FA fa20_15(.a(sum19[16]), .b(A[15] & B[20]), .ci(carry20[14]), .s(sum20[15]), .co(carry20[15]));
FA fa20_16(.a(sum19[17]), .b(A[16] & B[20]), .ci(carry20[15]), .s(sum20[16]), .co(carry20[16]));
FA fa20_17(.a(sum19[18]), .b(A[17] & B[20]), .ci(carry20[16]), .s(sum20[17]), .co(carry20[17]));
FA fa20_18(.a(sum19[19]), .b(A[18] & B[20]), .ci(carry20[17]), .s(sum20[18]), .co(carry20[18]));
FA fa20_19(.a(sum19[20]), .b(A[19] & B[20]), .ci(carry20[18]), .s(sum20[19]), .co(carry20[19]));
FA fa20_20(.a(sum19[21]), .b(A[20] & B[20]), .ci(carry20[19]), .s(sum20[20]), .co(carry20[20]));
FA fa20_21(.a(sum19[22]), .b(A[21] & B[20]), .ci(carry20[20]), .s(sum20[21]), .co(carry20[21]));
FA fa20_22(.a(sum19[23]), .b(A[22] & B[20]), .ci(carry20[21]), .s(sum20[22]), .co(carry20[22]));
FA fa20_23(.a(sum19[24]), .b(A[23] & B[20]), .ci(carry20[22]), .s(sum20[23]), .co(carry20[23]));
FA fa20_24(.a(sum19[25]), .b(A[24] & B[20]), .ci(carry20[23]), .s(sum20[24]), .co(carry20[24]));
FA fa20_25(.a(sum19[26]), .b(A[25] & B[20]), .ci(carry20[24]), .s(sum20[25]), .co(carry20[25]));
FA fa20_26(.a(sum19[27]), .b(A[26] & B[20]), .ci(carry20[25]), .s(sum20[26]), .co(carry20[26]));
FA fa20_27(.a(sum19[28]), .b(A[27] & B[20]), .ci(carry20[26]), .s(sum20[27]), .co(carry20[27]));
FA fa20_28(.a(sum19[29]), .b(A[28] & B[20]), .ci(carry20[27]), .s(sum20[28]), .co(carry20[28]));
FA fa20_29(.a(sum19[30]), .b(A[29] & B[20]), .ci(carry20[28]), .s(sum20[29]), .co(carry20[29]));
FA fa20_30(.a(sum19[31]), .b(A[30] & B[20]), .ci(carry20[29]), .s(sum20[30]), .co(carry20[30]));
FA fa20_31(.a(carry19[31]), .b(A[31] & B[20]), .ci(carry20[30]), .s(sum20[31]), .co(carry20[31]));
FA fa21_0(.a(sum20[1]), .b(A[0] & B[21]), .ci(1'b0), .s(Z[21]), .co(carry21[0]));
FA fa21_1(.a(sum20[2]), .b(A[1] & B[21]), .ci(carry21[0]), .s(sum21[1]), .co(carry21[1]));
FA fa21_2(.a(sum20[3]), .b(A[2] & B[21]), .ci(carry21[1]), .s(sum21[2]), .co(carry21[2]));
FA fa21_3(.a(sum20[4]), .b(A[3] & B[21]), .ci(carry21[2]), .s(sum21[3]), .co(carry21[3]));
FA fa21_4(.a(sum20[5]), .b(A[4] & B[21]), .ci(carry21[3]), .s(sum21[4]), .co(carry21[4]));
FA fa21_5(.a(sum20[6]), .b(A[5] & B[21]), .ci(carry21[4]), .s(sum21[5]), .co(carry21[5]));
FA fa21_6(.a(sum20[7]), .b(A[6] & B[21]), .ci(carry21[5]), .s(sum21[6]), .co(carry21[6]));
FA fa21_7(.a(sum20[8]), .b(A[7] & B[21]), .ci(carry21[6]), .s(sum21[7]), .co(carry21[7]));
FA fa21_8(.a(sum20[9]), .b(A[8] & B[21]), .ci(carry21[7]), .s(sum21[8]), .co(carry21[8]));
FA fa21_9(.a(sum20[10]), .b(A[9] & B[21]), .ci(carry21[8]), .s(sum21[9]), .co(carry21[9]));
FA fa21_10(.a(sum20[11]), .b(A[10] & B[21]), .ci(carry21[9]), .s(sum21[10]), .co(carry21[10]));
FA fa21_11(.a(sum20[12]), .b(A[11] & B[21]), .ci(carry21[10]), .s(sum21[11]), .co(carry21[11]));
FA fa21_12(.a(sum20[13]), .b(A[12] & B[21]), .ci(carry21[11]), .s(sum21[12]), .co(carry21[12]));
FA fa21_13(.a(sum20[14]), .b(A[13] & B[21]), .ci(carry21[12]), .s(sum21[13]), .co(carry21[13]));
FA fa21_14(.a(sum20[15]), .b(A[14] & B[21]), .ci(carry21[13]), .s(sum21[14]), .co(carry21[14]));
FA fa21_15(.a(sum20[16]), .b(A[15] & B[21]), .ci(carry21[14]), .s(sum21[15]), .co(carry21[15]));
FA fa21_16(.a(sum20[17]), .b(A[16] & B[21]), .ci(carry21[15]), .s(sum21[16]), .co(carry21[16]));
FA fa21_17(.a(sum20[18]), .b(A[17] & B[21]), .ci(carry21[16]), .s(sum21[17]), .co(carry21[17]));
FA fa21_18(.a(sum20[19]), .b(A[18] & B[21]), .ci(carry21[17]), .s(sum21[18]), .co(carry21[18]));
FA fa21_19(.a(sum20[20]), .b(A[19] & B[21]), .ci(carry21[18]), .s(sum21[19]), .co(carry21[19]));
FA fa21_20(.a(sum20[21]), .b(A[20] & B[21]), .ci(carry21[19]), .s(sum21[20]), .co(carry21[20]));
FA fa21_21(.a(sum20[22]), .b(A[21] & B[21]), .ci(carry21[20]), .s(sum21[21]), .co(carry21[21]));
FA fa21_22(.a(sum20[23]), .b(A[22] & B[21]), .ci(carry21[21]), .s(sum21[22]), .co(carry21[22]));
FA fa21_23(.a(sum20[24]), .b(A[23] & B[21]), .ci(carry21[22]), .s(sum21[23]), .co(carry21[23]));
FA fa21_24(.a(sum20[25]), .b(A[24] & B[21]), .ci(carry21[23]), .s(sum21[24]), .co(carry21[24]));
FA fa21_25(.a(sum20[26]), .b(A[25] & B[21]), .ci(carry21[24]), .s(sum21[25]), .co(carry21[25]));
FA fa21_26(.a(sum20[27]), .b(A[26] & B[21]), .ci(carry21[25]), .s(sum21[26]), .co(carry21[26]));
FA fa21_27(.a(sum20[28]), .b(A[27] & B[21]), .ci(carry21[26]), .s(sum21[27]), .co(carry21[27]));
FA fa21_28(.a(sum20[29]), .b(A[28] & B[21]), .ci(carry21[27]), .s(sum21[28]), .co(carry21[28]));
FA fa21_29(.a(sum20[30]), .b(A[29] & B[21]), .ci(carry21[28]), .s(sum21[29]), .co(carry21[29]));
FA fa21_30(.a(sum20[31]), .b(A[30] & B[21]), .ci(carry21[29]), .s(sum21[30]), .co(carry21[30]));
FA fa21_31(.a(carry20[31]), .b(A[31] & B[21]), .ci(carry21[30]), .s(sum21[31]), .co(carry21[31]));
FA fa22_0(.a(sum21[1]), .b(A[0] & B[22]), .ci(1'b0), .s(Z[22]), .co(carry22[0]));
FA fa22_1(.a(sum21[2]), .b(A[1] & B[22]), .ci(carry22[0]), .s(sum22[1]), .co(carry22[1]));
FA fa22_2(.a(sum21[3]), .b(A[2] & B[22]), .ci(carry22[1]), .s(sum22[2]), .co(carry22[2]));
FA fa22_3(.a(sum21[4]), .b(A[3] & B[22]), .ci(carry22[2]), .s(sum22[3]), .co(carry22[3]));
FA fa22_4(.a(sum21[5]), .b(A[4] & B[22]), .ci(carry22[3]), .s(sum22[4]), .co(carry22[4]));
FA fa22_5(.a(sum21[6]), .b(A[5] & B[22]), .ci(carry22[4]), .s(sum22[5]), .co(carry22[5]));
FA fa22_6(.a(sum21[7]), .b(A[6] & B[22]), .ci(carry22[5]), .s(sum22[6]), .co(carry22[6]));
FA fa22_7(.a(sum21[8]), .b(A[7] & B[22]), .ci(carry22[6]), .s(sum22[7]), .co(carry22[7]));
FA fa22_8(.a(sum21[9]), .b(A[8] & B[22]), .ci(carry22[7]), .s(sum22[8]), .co(carry22[8]));
FA fa22_9(.a(sum21[10]), .b(A[9] & B[22]), .ci(carry22[8]), .s(sum22[9]), .co(carry22[9]));
FA fa22_10(.a(sum21[11]), .b(A[10] & B[22]), .ci(carry22[9]), .s(sum22[10]), .co(carry22[10]));
FA fa22_11(.a(sum21[12]), .b(A[11] & B[22]), .ci(carry22[10]), .s(sum22[11]), .co(carry22[11]));
FA fa22_12(.a(sum21[13]), .b(A[12] & B[22]), .ci(carry22[11]), .s(sum22[12]), .co(carry22[12]));
FA fa22_13(.a(sum21[14]), .b(A[13] & B[22]), .ci(carry22[12]), .s(sum22[13]), .co(carry22[13]));
FA fa22_14(.a(sum21[15]), .b(A[14] & B[22]), .ci(carry22[13]), .s(sum22[14]), .co(carry22[14]));
FA fa22_15(.a(sum21[16]), .b(A[15] & B[22]), .ci(carry22[14]), .s(sum22[15]), .co(carry22[15]));
FA fa22_16(.a(sum21[17]), .b(A[16] & B[22]), .ci(carry22[15]), .s(sum22[16]), .co(carry22[16]));
FA fa22_17(.a(sum21[18]), .b(A[17] & B[22]), .ci(carry22[16]), .s(sum22[17]), .co(carry22[17]));
FA fa22_18(.a(sum21[19]), .b(A[18] & B[22]), .ci(carry22[17]), .s(sum22[18]), .co(carry22[18]));
FA fa22_19(.a(sum21[20]), .b(A[19] & B[22]), .ci(carry22[18]), .s(sum22[19]), .co(carry22[19]));
FA fa22_20(.a(sum21[21]), .b(A[20] & B[22]), .ci(carry22[19]), .s(sum22[20]), .co(carry22[20]));
FA fa22_21(.a(sum21[22]), .b(A[21] & B[22]), .ci(carry22[20]), .s(sum22[21]), .co(carry22[21]));
FA fa22_22(.a(sum21[23]), .b(A[22] & B[22]), .ci(carry22[21]), .s(sum22[22]), .co(carry22[22]));
FA fa22_23(.a(sum21[24]), .b(A[23] & B[22]), .ci(carry22[22]), .s(sum22[23]), .co(carry22[23]));
FA fa22_24(.a(sum21[25]), .b(A[24] & B[22]), .ci(carry22[23]), .s(sum22[24]), .co(carry22[24]));
FA fa22_25(.a(sum21[26]), .b(A[25] & B[22]), .ci(carry22[24]), .s(sum22[25]), .co(carry22[25]));
FA fa22_26(.a(sum21[27]), .b(A[26] & B[22]), .ci(carry22[25]), .s(sum22[26]), .co(carry22[26]));
FA fa22_27(.a(sum21[28]), .b(A[27] & B[22]), .ci(carry22[26]), .s(sum22[27]), .co(carry22[27]));
FA fa22_28(.a(sum21[29]), .b(A[28] & B[22]), .ci(carry22[27]), .s(sum22[28]), .co(carry22[28]));
FA fa22_29(.a(sum21[30]), .b(A[29] & B[22]), .ci(carry22[28]), .s(sum22[29]), .co(carry22[29]));
FA fa22_30(.a(sum21[31]), .b(A[30] & B[22]), .ci(carry22[29]), .s(sum22[30]), .co(carry22[30]));
FA fa22_31(.a(carry21[31]), .b(A[31] & B[22]), .ci(carry22[30]), .s(sum22[31]), .co(carry22[31]));
FA fa23_0(.a(sum22[1]), .b(A[0] & B[23]), .ci(1'b0), .s(Z[23]), .co(carry23[0]));
FA fa23_1(.a(sum22[2]), .b(A[1] & B[23]), .ci(carry23[0]), .s(sum23[1]), .co(carry23[1]));
FA fa23_2(.a(sum22[3]), .b(A[2] & B[23]), .ci(carry23[1]), .s(sum23[2]), .co(carry23[2]));
FA fa23_3(.a(sum22[4]), .b(A[3] & B[23]), .ci(carry23[2]), .s(sum23[3]), .co(carry23[3]));
FA fa23_4(.a(sum22[5]), .b(A[4] & B[23]), .ci(carry23[3]), .s(sum23[4]), .co(carry23[4]));
FA fa23_5(.a(sum22[6]), .b(A[5] & B[23]), .ci(carry23[4]), .s(sum23[5]), .co(carry23[5]));
FA fa23_6(.a(sum22[7]), .b(A[6] & B[23]), .ci(carry23[5]), .s(sum23[6]), .co(carry23[6]));
FA fa23_7(.a(sum22[8]), .b(A[7] & B[23]), .ci(carry23[6]), .s(sum23[7]), .co(carry23[7]));
FA fa23_8(.a(sum22[9]), .b(A[8] & B[23]), .ci(carry23[7]), .s(sum23[8]), .co(carry23[8]));
FA fa23_9(.a(sum22[10]), .b(A[9] & B[23]), .ci(carry23[8]), .s(sum23[9]), .co(carry23[9]));
FA fa23_10(.a(sum22[11]), .b(A[10] & B[23]), .ci(carry23[9]), .s(sum23[10]), .co(carry23[10]));
FA fa23_11(.a(sum22[12]), .b(A[11] & B[23]), .ci(carry23[10]), .s(sum23[11]), .co(carry23[11]));
FA fa23_12(.a(sum22[13]), .b(A[12] & B[23]), .ci(carry23[11]), .s(sum23[12]), .co(carry23[12]));
FA fa23_13(.a(sum22[14]), .b(A[13] & B[23]), .ci(carry23[12]), .s(sum23[13]), .co(carry23[13]));
FA fa23_14(.a(sum22[15]), .b(A[14] & B[23]), .ci(carry23[13]), .s(sum23[14]), .co(carry23[14]));
FA fa23_15(.a(sum22[16]), .b(A[15] & B[23]), .ci(carry23[14]), .s(sum23[15]), .co(carry23[15]));
FA fa23_16(.a(sum22[17]), .b(A[16] & B[23]), .ci(carry23[15]), .s(sum23[16]), .co(carry23[16]));
FA fa23_17(.a(sum22[18]), .b(A[17] & B[23]), .ci(carry23[16]), .s(sum23[17]), .co(carry23[17]));
FA fa23_18(.a(sum22[19]), .b(A[18] & B[23]), .ci(carry23[17]), .s(sum23[18]), .co(carry23[18]));
FA fa23_19(.a(sum22[20]), .b(A[19] & B[23]), .ci(carry23[18]), .s(sum23[19]), .co(carry23[19]));
FA fa23_20(.a(sum22[21]), .b(A[20] & B[23]), .ci(carry23[19]), .s(sum23[20]), .co(carry23[20]));
FA fa23_21(.a(sum22[22]), .b(A[21] & B[23]), .ci(carry23[20]), .s(sum23[21]), .co(carry23[21]));
FA fa23_22(.a(sum22[23]), .b(A[22] & B[23]), .ci(carry23[21]), .s(sum23[22]), .co(carry23[22]));
FA fa23_23(.a(sum22[24]), .b(A[23] & B[23]), .ci(carry23[22]), .s(sum23[23]), .co(carry23[23]));
FA fa23_24(.a(sum22[25]), .b(A[24] & B[23]), .ci(carry23[23]), .s(sum23[24]), .co(carry23[24]));
FA fa23_25(.a(sum22[26]), .b(A[25] & B[23]), .ci(carry23[24]), .s(sum23[25]), .co(carry23[25]));
FA fa23_26(.a(sum22[27]), .b(A[26] & B[23]), .ci(carry23[25]), .s(sum23[26]), .co(carry23[26]));
FA fa23_27(.a(sum22[28]), .b(A[27] & B[23]), .ci(carry23[26]), .s(sum23[27]), .co(carry23[27]));
FA fa23_28(.a(sum22[29]), .b(A[28] & B[23]), .ci(carry23[27]), .s(sum23[28]), .co(carry23[28]));
FA fa23_29(.a(sum22[30]), .b(A[29] & B[23]), .ci(carry23[28]), .s(sum23[29]), .co(carry23[29]));
FA fa23_30(.a(sum22[31]), .b(A[30] & B[23]), .ci(carry23[29]), .s(sum23[30]), .co(carry23[30]));
FA fa23_31(.a(carry22[31]), .b(A[31] & B[23]), .ci(carry23[30]), .s(sum23[31]), .co(carry23[31]));
FA fa24_0(.a(sum23[1]), .b(A[0] & B[24]), .ci(1'b0), .s(Z[24]), .co(carry24[0]));
FA fa24_1(.a(sum23[2]), .b(A[1] & B[24]), .ci(carry24[0]), .s(sum24[1]), .co(carry24[1]));
FA fa24_2(.a(sum23[3]), .b(A[2] & B[24]), .ci(carry24[1]), .s(sum24[2]), .co(carry24[2]));
FA fa24_3(.a(sum23[4]), .b(A[3] & B[24]), .ci(carry24[2]), .s(sum24[3]), .co(carry24[3]));
FA fa24_4(.a(sum23[5]), .b(A[4] & B[24]), .ci(carry24[3]), .s(sum24[4]), .co(carry24[4]));
FA fa24_5(.a(sum23[6]), .b(A[5] & B[24]), .ci(carry24[4]), .s(sum24[5]), .co(carry24[5]));
FA fa24_6(.a(sum23[7]), .b(A[6] & B[24]), .ci(carry24[5]), .s(sum24[6]), .co(carry24[6]));
FA fa24_7(.a(sum23[8]), .b(A[7] & B[24]), .ci(carry24[6]), .s(sum24[7]), .co(carry24[7]));
FA fa24_8(.a(sum23[9]), .b(A[8] & B[24]), .ci(carry24[7]), .s(sum24[8]), .co(carry24[8]));
FA fa24_9(.a(sum23[10]), .b(A[9] & B[24]), .ci(carry24[8]), .s(sum24[9]), .co(carry24[9]));
FA fa24_10(.a(sum23[11]), .b(A[10] & B[24]), .ci(carry24[9]), .s(sum24[10]), .co(carry24[10]));
FA fa24_11(.a(sum23[12]), .b(A[11] & B[24]), .ci(carry24[10]), .s(sum24[11]), .co(carry24[11]));
FA fa24_12(.a(sum23[13]), .b(A[12] & B[24]), .ci(carry24[11]), .s(sum24[12]), .co(carry24[12]));
FA fa24_13(.a(sum23[14]), .b(A[13] & B[24]), .ci(carry24[12]), .s(sum24[13]), .co(carry24[13]));
FA fa24_14(.a(sum23[15]), .b(A[14] & B[24]), .ci(carry24[13]), .s(sum24[14]), .co(carry24[14]));
FA fa24_15(.a(sum23[16]), .b(A[15] & B[24]), .ci(carry24[14]), .s(sum24[15]), .co(carry24[15]));
FA fa24_16(.a(sum23[17]), .b(A[16] & B[24]), .ci(carry24[15]), .s(sum24[16]), .co(carry24[16]));
FA fa24_17(.a(sum23[18]), .b(A[17] & B[24]), .ci(carry24[16]), .s(sum24[17]), .co(carry24[17]));
FA fa24_18(.a(sum23[19]), .b(A[18] & B[24]), .ci(carry24[17]), .s(sum24[18]), .co(carry24[18]));
FA fa24_19(.a(sum23[20]), .b(A[19] & B[24]), .ci(carry24[18]), .s(sum24[19]), .co(carry24[19]));
FA fa24_20(.a(sum23[21]), .b(A[20] & B[24]), .ci(carry24[19]), .s(sum24[20]), .co(carry24[20]));
FA fa24_21(.a(sum23[22]), .b(A[21] & B[24]), .ci(carry24[20]), .s(sum24[21]), .co(carry24[21]));
FA fa24_22(.a(sum23[23]), .b(A[22] & B[24]), .ci(carry24[21]), .s(sum24[22]), .co(carry24[22]));
FA fa24_23(.a(sum23[24]), .b(A[23] & B[24]), .ci(carry24[22]), .s(sum24[23]), .co(carry24[23]));
FA fa24_24(.a(sum23[25]), .b(A[24] & B[24]), .ci(carry24[23]), .s(sum24[24]), .co(carry24[24]));
FA fa24_25(.a(sum23[26]), .b(A[25] & B[24]), .ci(carry24[24]), .s(sum24[25]), .co(carry24[25]));
FA fa24_26(.a(sum23[27]), .b(A[26] & B[24]), .ci(carry24[25]), .s(sum24[26]), .co(carry24[26]));
FA fa24_27(.a(sum23[28]), .b(A[27] & B[24]), .ci(carry24[26]), .s(sum24[27]), .co(carry24[27]));
FA fa24_28(.a(sum23[29]), .b(A[28] & B[24]), .ci(carry24[27]), .s(sum24[28]), .co(carry24[28]));
FA fa24_29(.a(sum23[30]), .b(A[29] & B[24]), .ci(carry24[28]), .s(sum24[29]), .co(carry24[29]));
FA fa24_30(.a(sum23[31]), .b(A[30] & B[24]), .ci(carry24[29]), .s(sum24[30]), .co(carry24[30]));
FA fa24_31(.a(carry23[31]), .b(A[31] & B[24]), .ci(carry24[30]), .s(sum24[31]), .co(carry24[31]));
FA fa25_0(.a(sum24[1]), .b(A[0] & B[25]), .ci(1'b0), .s(Z[25]), .co(carry25[0]));
FA fa25_1(.a(sum24[2]), .b(A[1] & B[25]), .ci(carry25[0]), .s(sum25[1]), .co(carry25[1]));
FA fa25_2(.a(sum24[3]), .b(A[2] & B[25]), .ci(carry25[1]), .s(sum25[2]), .co(carry25[2]));
FA fa25_3(.a(sum24[4]), .b(A[3] & B[25]), .ci(carry25[2]), .s(sum25[3]), .co(carry25[3]));
FA fa25_4(.a(sum24[5]), .b(A[4] & B[25]), .ci(carry25[3]), .s(sum25[4]), .co(carry25[4]));
FA fa25_5(.a(sum24[6]), .b(A[5] & B[25]), .ci(carry25[4]), .s(sum25[5]), .co(carry25[5]));
FA fa25_6(.a(sum24[7]), .b(A[6] & B[25]), .ci(carry25[5]), .s(sum25[6]), .co(carry25[6]));
FA fa25_7(.a(sum24[8]), .b(A[7] & B[25]), .ci(carry25[6]), .s(sum25[7]), .co(carry25[7]));
FA fa25_8(.a(sum24[9]), .b(A[8] & B[25]), .ci(carry25[7]), .s(sum25[8]), .co(carry25[8]));
FA fa25_9(.a(sum24[10]), .b(A[9] & B[25]), .ci(carry25[8]), .s(sum25[9]), .co(carry25[9]));
FA fa25_10(.a(sum24[11]), .b(A[10] & B[25]), .ci(carry25[9]), .s(sum25[10]), .co(carry25[10]));
FA fa25_11(.a(sum24[12]), .b(A[11] & B[25]), .ci(carry25[10]), .s(sum25[11]), .co(carry25[11]));
FA fa25_12(.a(sum24[13]), .b(A[12] & B[25]), .ci(carry25[11]), .s(sum25[12]), .co(carry25[12]));
FA fa25_13(.a(sum24[14]), .b(A[13] & B[25]), .ci(carry25[12]), .s(sum25[13]), .co(carry25[13]));
FA fa25_14(.a(sum24[15]), .b(A[14] & B[25]), .ci(carry25[13]), .s(sum25[14]), .co(carry25[14]));
FA fa25_15(.a(sum24[16]), .b(A[15] & B[25]), .ci(carry25[14]), .s(sum25[15]), .co(carry25[15]));
FA fa25_16(.a(sum24[17]), .b(A[16] & B[25]), .ci(carry25[15]), .s(sum25[16]), .co(carry25[16]));
FA fa25_17(.a(sum24[18]), .b(A[17] & B[25]), .ci(carry25[16]), .s(sum25[17]), .co(carry25[17]));
FA fa25_18(.a(sum24[19]), .b(A[18] & B[25]), .ci(carry25[17]), .s(sum25[18]), .co(carry25[18]));
FA fa25_19(.a(sum24[20]), .b(A[19] & B[25]), .ci(carry25[18]), .s(sum25[19]), .co(carry25[19]));
FA fa25_20(.a(sum24[21]), .b(A[20] & B[25]), .ci(carry25[19]), .s(sum25[20]), .co(carry25[20]));
FA fa25_21(.a(sum24[22]), .b(A[21] & B[25]), .ci(carry25[20]), .s(sum25[21]), .co(carry25[21]));
FA fa25_22(.a(sum24[23]), .b(A[22] & B[25]), .ci(carry25[21]), .s(sum25[22]), .co(carry25[22]));
FA fa25_23(.a(sum24[24]), .b(A[23] & B[25]), .ci(carry25[22]), .s(sum25[23]), .co(carry25[23]));
FA fa25_24(.a(sum24[25]), .b(A[24] & B[25]), .ci(carry25[23]), .s(sum25[24]), .co(carry25[24]));
FA fa25_25(.a(sum24[26]), .b(A[25] & B[25]), .ci(carry25[24]), .s(sum25[25]), .co(carry25[25]));
FA fa25_26(.a(sum24[27]), .b(A[26] & B[25]), .ci(carry25[25]), .s(sum25[26]), .co(carry25[26]));
FA fa25_27(.a(sum24[28]), .b(A[27] & B[25]), .ci(carry25[26]), .s(sum25[27]), .co(carry25[27]));
FA fa25_28(.a(sum24[29]), .b(A[28] & B[25]), .ci(carry25[27]), .s(sum25[28]), .co(carry25[28]));
FA fa25_29(.a(sum24[30]), .b(A[29] & B[25]), .ci(carry25[28]), .s(sum25[29]), .co(carry25[29]));
FA fa25_30(.a(sum24[31]), .b(A[30] & B[25]), .ci(carry25[29]), .s(sum25[30]), .co(carry25[30]));
FA fa25_31(.a(carry24[31]), .b(A[31] & B[25]), .ci(carry25[30]), .s(sum25[31]), .co(carry25[31]));
FA fa26_0(.a(sum25[1]), .b(A[0] & B[26]), .ci(1'b0), .s(Z[26]), .co(carry26[0]));
FA fa26_1(.a(sum25[2]), .b(A[1] & B[26]), .ci(carry26[0]), .s(sum26[1]), .co(carry26[1]));
FA fa26_2(.a(sum25[3]), .b(A[2] & B[26]), .ci(carry26[1]), .s(sum26[2]), .co(carry26[2]));
FA fa26_3(.a(sum25[4]), .b(A[3] & B[26]), .ci(carry26[2]), .s(sum26[3]), .co(carry26[3]));
FA fa26_4(.a(sum25[5]), .b(A[4] & B[26]), .ci(carry26[3]), .s(sum26[4]), .co(carry26[4]));
FA fa26_5(.a(sum25[6]), .b(A[5] & B[26]), .ci(carry26[4]), .s(sum26[5]), .co(carry26[5]));
FA fa26_6(.a(sum25[7]), .b(A[6] & B[26]), .ci(carry26[5]), .s(sum26[6]), .co(carry26[6]));
FA fa26_7(.a(sum25[8]), .b(A[7] & B[26]), .ci(carry26[6]), .s(sum26[7]), .co(carry26[7]));
FA fa26_8(.a(sum25[9]), .b(A[8] & B[26]), .ci(carry26[7]), .s(sum26[8]), .co(carry26[8]));
FA fa26_9(.a(sum25[10]), .b(A[9] & B[26]), .ci(carry26[8]), .s(sum26[9]), .co(carry26[9]));
FA fa26_10(.a(sum25[11]), .b(A[10] & B[26]), .ci(carry26[9]), .s(sum26[10]), .co(carry26[10]));
FA fa26_11(.a(sum25[12]), .b(A[11] & B[26]), .ci(carry26[10]), .s(sum26[11]), .co(carry26[11]));
FA fa26_12(.a(sum25[13]), .b(A[12] & B[26]), .ci(carry26[11]), .s(sum26[12]), .co(carry26[12]));
FA fa26_13(.a(sum25[14]), .b(A[13] & B[26]), .ci(carry26[12]), .s(sum26[13]), .co(carry26[13]));
FA fa26_14(.a(sum25[15]), .b(A[14] & B[26]), .ci(carry26[13]), .s(sum26[14]), .co(carry26[14]));
FA fa26_15(.a(sum25[16]), .b(A[15] & B[26]), .ci(carry26[14]), .s(sum26[15]), .co(carry26[15]));
FA fa26_16(.a(sum25[17]), .b(A[16] & B[26]), .ci(carry26[15]), .s(sum26[16]), .co(carry26[16]));
FA fa26_17(.a(sum25[18]), .b(A[17] & B[26]), .ci(carry26[16]), .s(sum26[17]), .co(carry26[17]));
FA fa26_18(.a(sum25[19]), .b(A[18] & B[26]), .ci(carry26[17]), .s(sum26[18]), .co(carry26[18]));
FA fa26_19(.a(sum25[20]), .b(A[19] & B[26]), .ci(carry26[18]), .s(sum26[19]), .co(carry26[19]));
FA fa26_20(.a(sum25[21]), .b(A[20] & B[26]), .ci(carry26[19]), .s(sum26[20]), .co(carry26[20]));
FA fa26_21(.a(sum25[22]), .b(A[21] & B[26]), .ci(carry26[20]), .s(sum26[21]), .co(carry26[21]));
FA fa26_22(.a(sum25[23]), .b(A[22] & B[26]), .ci(carry26[21]), .s(sum26[22]), .co(carry26[22]));
FA fa26_23(.a(sum25[24]), .b(A[23] & B[26]), .ci(carry26[22]), .s(sum26[23]), .co(carry26[23]));
FA fa26_24(.a(sum25[25]), .b(A[24] & B[26]), .ci(carry26[23]), .s(sum26[24]), .co(carry26[24]));
FA fa26_25(.a(sum25[26]), .b(A[25] & B[26]), .ci(carry26[24]), .s(sum26[25]), .co(carry26[25]));
FA fa26_26(.a(sum25[27]), .b(A[26] & B[26]), .ci(carry26[25]), .s(sum26[26]), .co(carry26[26]));
FA fa26_27(.a(sum25[28]), .b(A[27] & B[26]), .ci(carry26[26]), .s(sum26[27]), .co(carry26[27]));
FA fa26_28(.a(sum25[29]), .b(A[28] & B[26]), .ci(carry26[27]), .s(sum26[28]), .co(carry26[28]));
FA fa26_29(.a(sum25[30]), .b(A[29] & B[26]), .ci(carry26[28]), .s(sum26[29]), .co(carry26[29]));
FA fa26_30(.a(sum25[31]), .b(A[30] & B[26]), .ci(carry26[29]), .s(sum26[30]), .co(carry26[30]));
FA fa26_31(.a(carry25[31]), .b(A[31] & B[26]), .ci(carry26[30]), .s(sum26[31]), .co(carry26[31]));
FA fa27_0(.a(sum26[1]), .b(A[0] & B[27]), .ci(1'b0), .s(Z[27]), .co(carry27[0]));
FA fa27_1(.a(sum26[2]), .b(A[1] & B[27]), .ci(carry27[0]), .s(sum27[1]), .co(carry27[1]));
FA fa27_2(.a(sum26[3]), .b(A[2] & B[27]), .ci(carry27[1]), .s(sum27[2]), .co(carry27[2]));
FA fa27_3(.a(sum26[4]), .b(A[3] & B[27]), .ci(carry27[2]), .s(sum27[3]), .co(carry27[3]));
FA fa27_4(.a(sum26[5]), .b(A[4] & B[27]), .ci(carry27[3]), .s(sum27[4]), .co(carry27[4]));
FA fa27_5(.a(sum26[6]), .b(A[5] & B[27]), .ci(carry27[4]), .s(sum27[5]), .co(carry27[5]));
FA fa27_6(.a(sum26[7]), .b(A[6] & B[27]), .ci(carry27[5]), .s(sum27[6]), .co(carry27[6]));
FA fa27_7(.a(sum26[8]), .b(A[7] & B[27]), .ci(carry27[6]), .s(sum27[7]), .co(carry27[7]));
FA fa27_8(.a(sum26[9]), .b(A[8] & B[27]), .ci(carry27[7]), .s(sum27[8]), .co(carry27[8]));
FA fa27_9(.a(sum26[10]), .b(A[9] & B[27]), .ci(carry27[8]), .s(sum27[9]), .co(carry27[9]));
FA fa27_10(.a(sum26[11]), .b(A[10] & B[27]), .ci(carry27[9]), .s(sum27[10]), .co(carry27[10]));
FA fa27_11(.a(sum26[12]), .b(A[11] & B[27]), .ci(carry27[10]), .s(sum27[11]), .co(carry27[11]));
FA fa27_12(.a(sum26[13]), .b(A[12] & B[27]), .ci(carry27[11]), .s(sum27[12]), .co(carry27[12]));
FA fa27_13(.a(sum26[14]), .b(A[13] & B[27]), .ci(carry27[12]), .s(sum27[13]), .co(carry27[13]));
FA fa27_14(.a(sum26[15]), .b(A[14] & B[27]), .ci(carry27[13]), .s(sum27[14]), .co(carry27[14]));
FA fa27_15(.a(sum26[16]), .b(A[15] & B[27]), .ci(carry27[14]), .s(sum27[15]), .co(carry27[15]));
FA fa27_16(.a(sum26[17]), .b(A[16] & B[27]), .ci(carry27[15]), .s(sum27[16]), .co(carry27[16]));
FA fa27_17(.a(sum26[18]), .b(A[17] & B[27]), .ci(carry27[16]), .s(sum27[17]), .co(carry27[17]));
FA fa27_18(.a(sum26[19]), .b(A[18] & B[27]), .ci(carry27[17]), .s(sum27[18]), .co(carry27[18]));
FA fa27_19(.a(sum26[20]), .b(A[19] & B[27]), .ci(carry27[18]), .s(sum27[19]), .co(carry27[19]));
FA fa27_20(.a(sum26[21]), .b(A[20] & B[27]), .ci(carry27[19]), .s(sum27[20]), .co(carry27[20]));
FA fa27_21(.a(sum26[22]), .b(A[21] & B[27]), .ci(carry27[20]), .s(sum27[21]), .co(carry27[21]));
FA fa27_22(.a(sum26[23]), .b(A[22] & B[27]), .ci(carry27[21]), .s(sum27[22]), .co(carry27[22]));
FA fa27_23(.a(sum26[24]), .b(A[23] & B[27]), .ci(carry27[22]), .s(sum27[23]), .co(carry27[23]));
FA fa27_24(.a(sum26[25]), .b(A[24] & B[27]), .ci(carry27[23]), .s(sum27[24]), .co(carry27[24]));
FA fa27_25(.a(sum26[26]), .b(A[25] & B[27]), .ci(carry27[24]), .s(sum27[25]), .co(carry27[25]));
FA fa27_26(.a(sum26[27]), .b(A[26] & B[27]), .ci(carry27[25]), .s(sum27[26]), .co(carry27[26]));
FA fa27_27(.a(sum26[28]), .b(A[27] & B[27]), .ci(carry27[26]), .s(sum27[27]), .co(carry27[27]));
FA fa27_28(.a(sum26[29]), .b(A[28] & B[27]), .ci(carry27[27]), .s(sum27[28]), .co(carry27[28]));
FA fa27_29(.a(sum26[30]), .b(A[29] & B[27]), .ci(carry27[28]), .s(sum27[29]), .co(carry27[29]));
FA fa27_30(.a(sum26[31]), .b(A[30] & B[27]), .ci(carry27[29]), .s(sum27[30]), .co(carry27[30]));
FA fa27_31(.a(carry26[31]), .b(A[31] & B[27]), .ci(carry27[30]), .s(sum27[31]), .co(carry27[31]));
FA fa28_0(.a(sum27[1]), .b(A[0] & B[28]), .ci(1'b0), .s(Z[28]), .co(carry28[0]));
FA fa28_1(.a(sum27[2]), .b(A[1] & B[28]), .ci(carry28[0]), .s(sum28[1]), .co(carry28[1]));
FA fa28_2(.a(sum27[3]), .b(A[2] & B[28]), .ci(carry28[1]), .s(sum28[2]), .co(carry28[2]));
FA fa28_3(.a(sum27[4]), .b(A[3] & B[28]), .ci(carry28[2]), .s(sum28[3]), .co(carry28[3]));
FA fa28_4(.a(sum27[5]), .b(A[4] & B[28]), .ci(carry28[3]), .s(sum28[4]), .co(carry28[4]));
FA fa28_5(.a(sum27[6]), .b(A[5] & B[28]), .ci(carry28[4]), .s(sum28[5]), .co(carry28[5]));
FA fa28_6(.a(sum27[7]), .b(A[6] & B[28]), .ci(carry28[5]), .s(sum28[6]), .co(carry28[6]));
FA fa28_7(.a(sum27[8]), .b(A[7] & B[28]), .ci(carry28[6]), .s(sum28[7]), .co(carry28[7]));
FA fa28_8(.a(sum27[9]), .b(A[8] & B[28]), .ci(carry28[7]), .s(sum28[8]), .co(carry28[8]));
FA fa28_9(.a(sum27[10]), .b(A[9] & B[28]), .ci(carry28[8]), .s(sum28[9]), .co(carry28[9]));
FA fa28_10(.a(sum27[11]), .b(A[10] & B[28]), .ci(carry28[9]), .s(sum28[10]), .co(carry28[10]));
FA fa28_11(.a(sum27[12]), .b(A[11] & B[28]), .ci(carry28[10]), .s(sum28[11]), .co(carry28[11]));
FA fa28_12(.a(sum27[13]), .b(A[12] & B[28]), .ci(carry28[11]), .s(sum28[12]), .co(carry28[12]));
FA fa28_13(.a(sum27[14]), .b(A[13] & B[28]), .ci(carry28[12]), .s(sum28[13]), .co(carry28[13]));
FA fa28_14(.a(sum27[15]), .b(A[14] & B[28]), .ci(carry28[13]), .s(sum28[14]), .co(carry28[14]));
FA fa28_15(.a(sum27[16]), .b(A[15] & B[28]), .ci(carry28[14]), .s(sum28[15]), .co(carry28[15]));
FA fa28_16(.a(sum27[17]), .b(A[16] & B[28]), .ci(carry28[15]), .s(sum28[16]), .co(carry28[16]));
FA fa28_17(.a(sum27[18]), .b(A[17] & B[28]), .ci(carry28[16]), .s(sum28[17]), .co(carry28[17]));
FA fa28_18(.a(sum27[19]), .b(A[18] & B[28]), .ci(carry28[17]), .s(sum28[18]), .co(carry28[18]));
FA fa28_19(.a(sum27[20]), .b(A[19] & B[28]), .ci(carry28[18]), .s(sum28[19]), .co(carry28[19]));
FA fa28_20(.a(sum27[21]), .b(A[20] & B[28]), .ci(carry28[19]), .s(sum28[20]), .co(carry28[20]));
FA fa28_21(.a(sum27[22]), .b(A[21] & B[28]), .ci(carry28[20]), .s(sum28[21]), .co(carry28[21]));
FA fa28_22(.a(sum27[23]), .b(A[22] & B[28]), .ci(carry28[21]), .s(sum28[22]), .co(carry28[22]));
FA fa28_23(.a(sum27[24]), .b(A[23] & B[28]), .ci(carry28[22]), .s(sum28[23]), .co(carry28[23]));
FA fa28_24(.a(sum27[25]), .b(A[24] & B[28]), .ci(carry28[23]), .s(sum28[24]), .co(carry28[24]));
FA fa28_25(.a(sum27[26]), .b(A[25] & B[28]), .ci(carry28[24]), .s(sum28[25]), .co(carry28[25]));
FA fa28_26(.a(sum27[27]), .b(A[26] & B[28]), .ci(carry28[25]), .s(sum28[26]), .co(carry28[26]));
FA fa28_27(.a(sum27[28]), .b(A[27] & B[28]), .ci(carry28[26]), .s(sum28[27]), .co(carry28[27]));
FA fa28_28(.a(sum27[29]), .b(A[28] & B[28]), .ci(carry28[27]), .s(sum28[28]), .co(carry28[28]));
FA fa28_29(.a(sum27[30]), .b(A[29] & B[28]), .ci(carry28[28]), .s(sum28[29]), .co(carry28[29]));
FA fa28_30(.a(sum27[31]), .b(A[30] & B[28]), .ci(carry28[29]), .s(sum28[30]), .co(carry28[30]));
FA fa28_31(.a(carry27[31]), .b(A[31] & B[28]), .ci(carry28[30]), .s(sum28[31]), .co(carry28[31]));
FA fa29_0(.a(sum28[1]), .b(A[0] & B[29]), .ci(1'b0), .s(Z[29]), .co(carry29[0]));
FA fa29_1(.a(sum28[2]), .b(A[1] & B[29]), .ci(carry29[0]), .s(sum29[1]), .co(carry29[1]));
FA fa29_2(.a(sum28[3]), .b(A[2] & B[29]), .ci(carry29[1]), .s(sum29[2]), .co(carry29[2]));
FA fa29_3(.a(sum28[4]), .b(A[3] & B[29]), .ci(carry29[2]), .s(sum29[3]), .co(carry29[3]));
FA fa29_4(.a(sum28[5]), .b(A[4] & B[29]), .ci(carry29[3]), .s(sum29[4]), .co(carry29[4]));
FA fa29_5(.a(sum28[6]), .b(A[5] & B[29]), .ci(carry29[4]), .s(sum29[5]), .co(carry29[5]));
FA fa29_6(.a(sum28[7]), .b(A[6] & B[29]), .ci(carry29[5]), .s(sum29[6]), .co(carry29[6]));
FA fa29_7(.a(sum28[8]), .b(A[7] & B[29]), .ci(carry29[6]), .s(sum29[7]), .co(carry29[7]));
FA fa29_8(.a(sum28[9]), .b(A[8] & B[29]), .ci(carry29[7]), .s(sum29[8]), .co(carry29[8]));
FA fa29_9(.a(sum28[10]), .b(A[9] & B[29]), .ci(carry29[8]), .s(sum29[9]), .co(carry29[9]));
FA fa29_10(.a(sum28[11]), .b(A[10] & B[29]), .ci(carry29[9]), .s(sum29[10]), .co(carry29[10]));
FA fa29_11(.a(sum28[12]), .b(A[11] & B[29]), .ci(carry29[10]), .s(sum29[11]), .co(carry29[11]));
FA fa29_12(.a(sum28[13]), .b(A[12] & B[29]), .ci(carry29[11]), .s(sum29[12]), .co(carry29[12]));
FA fa29_13(.a(sum28[14]), .b(A[13] & B[29]), .ci(carry29[12]), .s(sum29[13]), .co(carry29[13]));
FA fa29_14(.a(sum28[15]), .b(A[14] & B[29]), .ci(carry29[13]), .s(sum29[14]), .co(carry29[14]));
FA fa29_15(.a(sum28[16]), .b(A[15] & B[29]), .ci(carry29[14]), .s(sum29[15]), .co(carry29[15]));
FA fa29_16(.a(sum28[17]), .b(A[16] & B[29]), .ci(carry29[15]), .s(sum29[16]), .co(carry29[16]));
FA fa29_17(.a(sum28[18]), .b(A[17] & B[29]), .ci(carry29[16]), .s(sum29[17]), .co(carry29[17]));
FA fa29_18(.a(sum28[19]), .b(A[18] & B[29]), .ci(carry29[17]), .s(sum29[18]), .co(carry29[18]));
FA fa29_19(.a(sum28[20]), .b(A[19] & B[29]), .ci(carry29[18]), .s(sum29[19]), .co(carry29[19]));
FA fa29_20(.a(sum28[21]), .b(A[20] & B[29]), .ci(carry29[19]), .s(sum29[20]), .co(carry29[20]));
FA fa29_21(.a(sum28[22]), .b(A[21] & B[29]), .ci(carry29[20]), .s(sum29[21]), .co(carry29[21]));
FA fa29_22(.a(sum28[23]), .b(A[22] & B[29]), .ci(carry29[21]), .s(sum29[22]), .co(carry29[22]));
FA fa29_23(.a(sum28[24]), .b(A[23] & B[29]), .ci(carry29[22]), .s(sum29[23]), .co(carry29[23]));
FA fa29_24(.a(sum28[25]), .b(A[24] & B[29]), .ci(carry29[23]), .s(sum29[24]), .co(carry29[24]));
FA fa29_25(.a(sum28[26]), .b(A[25] & B[29]), .ci(carry29[24]), .s(sum29[25]), .co(carry29[25]));
FA fa29_26(.a(sum28[27]), .b(A[26] & B[29]), .ci(carry29[25]), .s(sum29[26]), .co(carry29[26]));
FA fa29_27(.a(sum28[28]), .b(A[27] & B[29]), .ci(carry29[26]), .s(sum29[27]), .co(carry29[27]));
FA fa29_28(.a(sum28[29]), .b(A[28] & B[29]), .ci(carry29[27]), .s(sum29[28]), .co(carry29[28]));
FA fa29_29(.a(sum28[30]), .b(A[29] & B[29]), .ci(carry29[28]), .s(sum29[29]), .co(carry29[29]));
FA fa29_30(.a(sum28[31]), .b(A[30] & B[29]), .ci(carry29[29]), .s(sum29[30]), .co(carry29[30]));
FA fa29_31(.a(carry28[31]), .b(A[31] & B[29]), .ci(carry29[30]), .s(sum29[31]), .co(carry29[31]));
FA fa30_0(.a(sum29[1]), .b(A[0] & B[30]), .ci(1'b0), .s(Z[30]), .co(carry30[0]));
FA fa30_1(.a(sum29[2]), .b(A[1] & B[30]), .ci(carry30[0]), .s(sum30[1]), .co(carry30[1]));
FA fa30_2(.a(sum29[3]), .b(A[2] & B[30]), .ci(carry30[1]), .s(sum30[2]), .co(carry30[2]));
FA fa30_3(.a(sum29[4]), .b(A[3] & B[30]), .ci(carry30[2]), .s(sum30[3]), .co(carry30[3]));
FA fa30_4(.a(sum29[5]), .b(A[4] & B[30]), .ci(carry30[3]), .s(sum30[4]), .co(carry30[4]));
FA fa30_5(.a(sum29[6]), .b(A[5] & B[30]), .ci(carry30[4]), .s(sum30[5]), .co(carry30[5]));
FA fa30_6(.a(sum29[7]), .b(A[6] & B[30]), .ci(carry30[5]), .s(sum30[6]), .co(carry30[6]));
FA fa30_7(.a(sum29[8]), .b(A[7] & B[30]), .ci(carry30[6]), .s(sum30[7]), .co(carry30[7]));
FA fa30_8(.a(sum29[9]), .b(A[8] & B[30]), .ci(carry30[7]), .s(sum30[8]), .co(carry30[8]));
FA fa30_9(.a(sum29[10]), .b(A[9] & B[30]), .ci(carry30[8]), .s(sum30[9]), .co(carry30[9]));
FA fa30_10(.a(sum29[11]), .b(A[10] & B[30]), .ci(carry30[9]), .s(sum30[10]), .co(carry30[10]));
FA fa30_11(.a(sum29[12]), .b(A[11] & B[30]), .ci(carry30[10]), .s(sum30[11]), .co(carry30[11]));
FA fa30_12(.a(sum29[13]), .b(A[12] & B[30]), .ci(carry30[11]), .s(sum30[12]), .co(carry30[12]));
FA fa30_13(.a(sum29[14]), .b(A[13] & B[30]), .ci(carry30[12]), .s(sum30[13]), .co(carry30[13]));
FA fa30_14(.a(sum29[15]), .b(A[14] & B[30]), .ci(carry30[13]), .s(sum30[14]), .co(carry30[14]));
FA fa30_15(.a(sum29[16]), .b(A[15] & B[30]), .ci(carry30[14]), .s(sum30[15]), .co(carry30[15]));
FA fa30_16(.a(sum29[17]), .b(A[16] & B[30]), .ci(carry30[15]), .s(sum30[16]), .co(carry30[16]));
FA fa30_17(.a(sum29[18]), .b(A[17] & B[30]), .ci(carry30[16]), .s(sum30[17]), .co(carry30[17]));
FA fa30_18(.a(sum29[19]), .b(A[18] & B[30]), .ci(carry30[17]), .s(sum30[18]), .co(carry30[18]));
FA fa30_19(.a(sum29[20]), .b(A[19] & B[30]), .ci(carry30[18]), .s(sum30[19]), .co(carry30[19]));
FA fa30_20(.a(sum29[21]), .b(A[20] & B[30]), .ci(carry30[19]), .s(sum30[20]), .co(carry30[20]));
FA fa30_21(.a(sum29[22]), .b(A[21] & B[30]), .ci(carry30[20]), .s(sum30[21]), .co(carry30[21]));
FA fa30_22(.a(sum29[23]), .b(A[22] & B[30]), .ci(carry30[21]), .s(sum30[22]), .co(carry30[22]));
FA fa30_23(.a(sum29[24]), .b(A[23] & B[30]), .ci(carry30[22]), .s(sum30[23]), .co(carry30[23]));
FA fa30_24(.a(sum29[25]), .b(A[24] & B[30]), .ci(carry30[23]), .s(sum30[24]), .co(carry30[24]));
FA fa30_25(.a(sum29[26]), .b(A[25] & B[30]), .ci(carry30[24]), .s(sum30[25]), .co(carry30[25]));
FA fa30_26(.a(sum29[27]), .b(A[26] & B[30]), .ci(carry30[25]), .s(sum30[26]), .co(carry30[26]));
FA fa30_27(.a(sum29[28]), .b(A[27] & B[30]), .ci(carry30[26]), .s(sum30[27]), .co(carry30[27]));
FA fa30_28(.a(sum29[29]), .b(A[28] & B[30]), .ci(carry30[27]), .s(sum30[28]), .co(carry30[28]));
FA fa30_29(.a(sum29[30]), .b(A[29] & B[30]), .ci(carry30[28]), .s(sum30[29]), .co(carry30[29]));
FA fa30_30(.a(sum29[31]), .b(A[30] & B[30]), .ci(carry30[29]), .s(sum30[30]), .co(carry30[30]));
FA fa30_31(.a(carry29[31]), .b(A[31] & B[30]), .ci(carry30[30]), .s(sum30[31]), .co(carry30[31]));
FA fa31_0(.a(sum30[1]), .b(A[0] & B[31]), .ci(1'b0), .s(Z[31]), .co(carry31[0]));
FA fa31_1(.a(sum30[2]), .b(A[1] & B[31]), .ci(carry31[0]), .s(sum31[1]), .co(carry31[1]));
FA fa31_2(.a(sum30[3]), .b(A[2] & B[31]), .ci(carry31[1]), .s(sum31[2]), .co(carry31[2]));
FA fa31_3(.a(sum30[4]), .b(A[3] & B[31]), .ci(carry31[2]), .s(sum31[3]), .co(carry31[3]));
FA fa31_4(.a(sum30[5]), .b(A[4] & B[31]), .ci(carry31[3]), .s(sum31[4]), .co(carry31[4]));
FA fa31_5(.a(sum30[6]), .b(A[5] & B[31]), .ci(carry31[4]), .s(sum31[5]), .co(carry31[5]));
FA fa31_6(.a(sum30[7]), .b(A[6] & B[31]), .ci(carry31[5]), .s(sum31[6]), .co(carry31[6]));
FA fa31_7(.a(sum30[8]), .b(A[7] & B[31]), .ci(carry31[6]), .s(sum31[7]), .co(carry31[7]));
FA fa31_8(.a(sum30[9]), .b(A[8] & B[31]), .ci(carry31[7]), .s(sum31[8]), .co(carry31[8]));
FA fa31_9(.a(sum30[10]), .b(A[9] & B[31]), .ci(carry31[8]), .s(sum31[9]), .co(carry31[9]));
FA fa31_10(.a(sum30[11]), .b(A[10] & B[31]), .ci(carry31[9]), .s(sum31[10]), .co(carry31[10]));
FA fa31_11(.a(sum30[12]), .b(A[11] & B[31]), .ci(carry31[10]), .s(sum31[11]), .co(carry31[11]));
FA fa31_12(.a(sum30[13]), .b(A[12] & B[31]), .ci(carry31[11]), .s(sum31[12]), .co(carry31[12]));
FA fa31_13(.a(sum30[14]), .b(A[13] & B[31]), .ci(carry31[12]), .s(sum31[13]), .co(carry31[13]));
FA fa31_14(.a(sum30[15]), .b(A[14] & B[31]), .ci(carry31[13]), .s(sum31[14]), .co(carry31[14]));
FA fa31_15(.a(sum30[16]), .b(A[15] & B[31]), .ci(carry31[14]), .s(sum31[15]), .co(carry31[15]));
FA fa31_16(.a(sum30[17]), .b(A[16] & B[31]), .ci(carry31[15]), .s(sum31[16]), .co(carry31[16]));
FA fa31_17(.a(sum30[18]), .b(A[17] & B[31]), .ci(carry31[16]), .s(sum31[17]), .co(carry31[17]));
FA fa31_18(.a(sum30[19]), .b(A[18] & B[31]), .ci(carry31[17]), .s(sum31[18]), .co(carry31[18]));
FA fa31_19(.a(sum30[20]), .b(A[19] & B[31]), .ci(carry31[18]), .s(sum31[19]), .co(carry31[19]));
FA fa31_20(.a(sum30[21]), .b(A[20] & B[31]), .ci(carry31[19]), .s(sum31[20]), .co(carry31[20]));
FA fa31_21(.a(sum30[22]), .b(A[21] & B[31]), .ci(carry31[20]), .s(sum31[21]), .co(carry31[21]));
FA fa31_22(.a(sum30[23]), .b(A[22] & B[31]), .ci(carry31[21]), .s(sum31[22]), .co(carry31[22]));
FA fa31_23(.a(sum30[24]), .b(A[23] & B[31]), .ci(carry31[22]), .s(sum31[23]), .co(carry31[23]));
FA fa31_24(.a(sum30[25]), .b(A[24] & B[31]), .ci(carry31[23]), .s(sum31[24]), .co(carry31[24]));
FA fa31_25(.a(sum30[26]), .b(A[25] & B[31]), .ci(carry31[24]), .s(sum31[25]), .co(carry31[25]));
FA fa31_26(.a(sum30[27]), .b(A[26] & B[31]), .ci(carry31[25]), .s(sum31[26]), .co(carry31[26]));
FA fa31_27(.a(sum30[28]), .b(A[27] & B[31]), .ci(carry31[26]), .s(sum31[27]), .co(carry31[27]));
FA fa31_28(.a(sum30[29]), .b(A[28] & B[31]), .ci(carry31[27]), .s(sum31[28]), .co(carry31[28]));
FA fa31_29(.a(sum30[30]), .b(A[29] & B[31]), .ci(carry31[28]), .s(sum31[29]), .co(carry31[29]));
FA fa31_30(.a(sum30[31]), .b(A[30] & B[31]), .ci(carry31[29]), .s(sum31[30]), .co(carry31[30]));
FA fa31_31(.a(carry30[31]), .b(A[31] & B[31]), .ci(carry31[30]), .s(sum31[31]), .co(carry31[31]));

assign Z[0] = sum0[0];
assign Z[1] = sum1[0];
assign Z[2] = sum2[0];
assign Z[3] = sum3[0];
assign Z[4] = sum4[0];
assign Z[5] = sum5[0];
assign Z[6] = sum6[0];
assign Z[7] = sum7[0];
assign Z[8] = sum8[0];
assign Z[9] = sum9[0];
assign Z[10] = sum10[0];
assign Z[11] = sum11[0];
assign Z[12] = sum12[0];
assign Z[13] = sum13[0];
assign Z[14] = sum14[0];
assign Z[15] = sum15[0];
assign Z[16] = sum16[0];
assign Z[17] = sum17[0];
assign Z[18] = sum18[0];
assign Z[19] = sum19[0];
assign Z[20] = sum20[0];
assign Z[21] = sum21[0];
assign Z[22] = sum22[0];
assign Z[23] = sum23[0];
assign Z[24] = sum24[0];
assign Z[25] = sum25[0];
assign Z[26] = sum26[0];
assign Z[27] = sum27[0];
assign Z[28] = sum28[0];
assign Z[29] = sum29[0];
assign Z[30] = sum30[0];
assign Z[62:31] = sum31;
assign Z[63] = carry31[31];


endmodule